// 6502 Final Netlist with CTS and ECO
// Design cells: 28819
// CTS/ECO cells: 0
// Total: 28819

module 6502_final (clk, rst_n, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, in_38, in_39, oeb_0, oeb_1, oeb_2, oeb_3, oeb_4, oeb_5, oeb_6, oeb_7, oeb_8, oeb_9, oeb_10, oeb_11, oeb_12, oeb_13, oeb_14, oeb_15, oeb_16, oeb_17, oeb_18, oeb_19, oeb_20, oeb_21, oeb_22, oeb_23, oeb_24, oeb_25, oeb_26, oeb_27, oeb_28, oeb_29, oeb_30, oeb_31, oeb_32, oeb_33, oeb_34, oeb_35, oeb_36, oeb_37, oeb_38, oeb_39, out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21, out_22, out_23, out_24, out_25, out_26, out_27, out_28, out_29, out_30, out_31, out_32, out_33, out_34, out_35, out_36, out_37, out_38, out_39);

  input clk;
  input rst_n;
  input in_0;
  input in_1;
  input in_2;
  input in_3;
  input in_4;
  input in_5;
  input in_6;
  input in_7;
  input in_8;
  input in_9;
  input in_10;
  input in_11;
  input in_12;
  input in_13;
  input in_14;
  input in_15;
  input in_16;
  input in_17;
  input in_18;
  input in_19;
  input in_20;
  input in_21;
  input in_22;
  input in_23;
  input in_24;
  input in_25;
  input in_26;
  input in_27;
  input in_28;
  input in_29;
  input in_30;
  input in_31;
  input in_32;
  input in_33;
  input in_34;
  input in_35;
  input in_36;
  input in_37;
  input in_38;
  input in_39;
  output oeb_0;
  output oeb_1;
  output oeb_2;
  output oeb_3;
  output oeb_4;
  output oeb_5;
  output oeb_6;
  output oeb_7;
  output oeb_8;
  output oeb_9;
  output oeb_10;
  output oeb_11;
  output oeb_12;
  output oeb_13;
  output oeb_14;
  output oeb_15;
  output oeb_16;
  output oeb_17;
  output oeb_18;
  output oeb_19;
  output oeb_20;
  output oeb_21;
  output oeb_22;
  output oeb_23;
  output oeb_24;
  output oeb_25;
  output oeb_26;
  output oeb_27;
  output oeb_28;
  output oeb_29;
  output oeb_30;
  output oeb_31;
  output oeb_32;
  output oeb_33;
  output oeb_34;
  output oeb_35;
  output oeb_36;
  output oeb_37;
  output oeb_38;
  output oeb_39;
  output out_0;
  output out_1;
  output out_2;
  output out_3;
  output out_4;
  output out_5;
  output out_6;
  output out_7;
  output out_8;
  output out_9;
  output out_10;
  output out_11;
  output out_12;
  output out_13;
  output out_14;
  output out_15;
  output out_16;
  output out_17;
  output out_18;
  output out_19;
  output out_20;
  output out_21;
  output out_22;
  output out_23;
  output out_24;
  output out_25;
  output out_26;
  output out_27;
  output out_28;
  output out_29;
  output out_30;
  output out_31;
  output out_32;
  output out_33;
  output out_34;
  output out_35;
  output out_36;
  output out_37;
  output out_38;
  output out_39;

  // Internal nets
  wire 100;
  wire 1000;
  wire 1001;
  wire 1002;
  wire 1003;
  wire 1004;
  wire 1005;
  wire 1006;
  wire 1007;
  wire 1008;
  wire 1009;
  wire 101;
  wire 1010;
  wire 1011;
  wire 1012;
  wire 1013;
  wire 1014;
  wire 1015;
  wire 1016;
  wire 1017;
  wire 1018;
  wire 1019;
  wire 102;
  wire 1020;
  wire 1021;
  wire 1022;
  wire 1023;
  wire 1024;
  wire 1025;
  wire 1026;
  wire 1027;
  wire 1028;
  wire 1029;
  wire 103;
  wire 1030;
  wire 1031;
  wire 1032;
  wire 1033;
  wire 1034;
  wire 1035;
  wire 1036;
  wire 1037;
  wire 1038;
  wire 1039;
  wire 104;
  wire 1040;
  wire 1041;
  wire 1042;
  wire 1043;
  wire 1044;
  wire 1045;
  wire 1046;
  wire 1047;
  wire 1048;
  wire 1049;
  wire 105;
  wire 1050;
  wire 1051;
  wire 1052;
  wire 1053;
  wire 1054;
  wire 1055;
  wire 1056;
  wire 1057;
  wire 1058;
  wire 1059;
  wire 106;
  wire 1060;
  wire 1061;
  wire 1062;
  wire 1063;
  wire 1064;
  wire 1065;
  wire 1066;
  wire 1067;
  wire 1068;
  wire 1069;
  wire 107;
  wire 1070;
  wire 1071;
  wire 1072;
  wire 1073;
  wire 1074;
  wire 1075;
  wire 1076;
  wire 1077;
  wire 1078;
  wire 1079;
  wire 108;
  wire 1080;
  wire 1081;
  wire 1082;
  wire 1083;
  wire 1084;
  wire 1085;
  wire 1086;
  wire 1087;
  wire 1088;
  wire 1089;
  wire 109;
  wire 1090;
  wire 1091;
  wire 1092;
  wire 1093;
  wire 1094;
  wire 1095;
  wire 1096;
  wire 1097;
  wire 1098;
  wire 1099;
  wire 110;
  wire 1100;
  wire 1101;
  wire 1102;
  wire 1103;
  wire 1104;
  wire 1105;
  wire 1106;
  wire 1107;
  wire 1108;
  wire 1109;
  wire 111;
  wire 1110;
  wire 1111;
  wire 1112;
  wire 1113;
  wire 1114;
  wire 1115;
  wire 1116;
  wire 1117;
  wire 1118;
  wire 1119;
  wire 112;
  wire 1120;
  wire 1121;
  wire 1122;
  wire 1123;
  wire 1124;
  wire 1125;
  wire 1126;
  wire 1127;
  wire 1128;
  wire 1129;
  wire 113;
  wire 1130;
  wire 1131;
  wire 1132;
  wire 1133;
  wire 1134;
  wire 1135;
  wire 1136;
  wire 1137;
  wire 1138;
  wire 1139;
  wire 114;
  wire 1140;
  wire 1141;
  wire 1142;
  wire 1143;
  wire 1144;
  wire 1145;
  wire 1146;
  wire 1147;
  wire 1148;
  wire 1149;
  wire 115;
  wire 1150;
  wire 1151;
  wire 1152;
  wire 1153;
  wire 1154;
  wire 1155;
  wire 1156;
  wire 1157;
  wire 1158;
  wire 1159;
  wire 116;
  wire 1160;
  wire 1161;
  wire 1162;
  wire 1163;
  wire 1164;
  wire 1165;
  wire 1166;
  wire 1167;
  wire 1168;
  wire 1169;
  wire 117;
  wire 1170;
  wire 1171;
  wire 1172;
  wire 1173;
  wire 1174;
  wire 1175;
  wire 1176;
  wire 1177;
  wire 1178;
  wire 1179;
  wire 118;
  wire 1180;
  wire 1181;
  wire 1182;
  wire 1183;
  wire 1184;
  wire 1185;
  wire 1186;
  wire 1187;
  wire 1188;
  wire 1189;
  wire 119;
  wire 1190;
  wire 1191;
  wire 1192;
  wire 1193;
  wire 1194;
  wire 1195;
  wire 1196;
  wire 1197;
  wire 1198;
  wire 1199;
  wire 120;
  wire 1200;
  wire 1201;
  wire 1202;
  wire 1203;
  wire 1204;
  wire 1205;
  wire 1206;
  wire 1207;
  wire 1208;
  wire 1209;
  wire 121;
  wire 1210;
  wire 1211;
  wire 1212;
  wire 1213;
  wire 1214;
  wire 1215;
  wire 1216;
  wire 1217;
  wire 1218;
  wire 1219;
  wire 122;
  wire 1220;
  wire 1221;
  wire 1222;
  wire 1223;
  wire 1224;
  wire 1225;
  wire 1226;
  wire 1227;
  wire 1228;
  wire 1229;
  wire 123;
  wire 1230;
  wire 1231;
  wire 1232;
  wire 1233;
  wire 1234;
  wire 1235;
  wire 1236;
  wire 1237;
  wire 1238;
  wire 1239;
  wire 124;
  wire 1240;
  wire 1241;
  wire 1242;
  wire 1243;
  wire 1244;
  wire 1245;
  wire 1246;
  wire 1247;
  wire 1248;
  wire 1249;
  wire 125;
  wire 1250;
  wire 1251;
  wire 1252;
  wire 1253;
  wire 1254;
  wire 1255;
  wire 1256;
  wire 1257;
  wire 1258;
  wire 1259;
  wire 126;
  wire 1260;
  wire 1261;
  wire 1262;
  wire 1263;
  wire 1264;
  wire 1265;
  wire 1266;
  wire 1267;
  wire 1268;
  wire 1269;
  wire 127;
  wire 1270;
  wire 1271;
  wire 1272;
  wire 1273;
  wire 1274;
  wire 1275;
  wire 1276;
  wire 1277;
  wire 1278;
  wire 1279;
  wire 128;
  wire 1280;
  wire 1281;
  wire 1282;
  wire 1283;
  wire 1284;
  wire 1285;
  wire 1286;
  wire 1287;
  wire 1288;
  wire 1289;
  wire 129;
  wire 1290;
  wire 1291;
  wire 1292;
  wire 1293;
  wire 1294;
  wire 1295;
  wire 1296;
  wire 1297;
  wire 1298;
  wire 1299;
  wire 130;
  wire 1300;
  wire 1301;
  wire 1302;
  wire 1303;
  wire 1304;
  wire 1305;
  wire 1306;
  wire 1307;
  wire 1308;
  wire 1309;
  wire 131;
  wire 1310;
  wire 1311;
  wire 1312;
  wire 1313;
  wire 1314;
  wire 1315;
  wire 1316;
  wire 1317;
  wire 1318;
  wire 1319;
  wire 132;
  wire 1320;
  wire 1321;
  wire 1322;
  wire 1323;
  wire 1324;
  wire 1325;
  wire 1326;
  wire 1327;
  wire 1328;
  wire 1329;
  wire 133;
  wire 1330;
  wire 1331;
  wire 1332;
  wire 1333;
  wire 1334;
  wire 1335;
  wire 1336;
  wire 1337;
  wire 1338;
  wire 1339;
  wire 134;
  wire 1340;
  wire 1341;
  wire 1342;
  wire 1343;
  wire 1344;
  wire 1345;
  wire 1346;
  wire 1347;
  wire 1348;
  wire 1349;
  wire 135;
  wire 1350;
  wire 1351;
  wire 1352;
  wire 1353;
  wire 1354;
  wire 1355;
  wire 1356;
  wire 1357;
  wire 1358;
  wire 1359;
  wire 136;
  wire 1360;
  wire 1361;
  wire 1362;
  wire 1363;
  wire 1364;
  wire 1365;
  wire 1366;
  wire 1367;
  wire 1368;
  wire 1369;
  wire 137;
  wire 1370;
  wire 1371;
  wire 1372;
  wire 1373;
  wire 1374;
  wire 1375;
  wire 1376;
  wire 1377;
  wire 1378;
  wire 1379;
  wire 138;
  wire 1380;
  wire 1381;
  wire 1382;
  wire 1383;
  wire 1384;
  wire 1385;
  wire 1386;
  wire 1387;
  wire 1388;
  wire 1389;
  wire 139;
  wire 1390;
  wire 1391;
  wire 1392;
  wire 1393;
  wire 1394;
  wire 1395;
  wire 1396;
  wire 1397;
  wire 1398;
  wire 1399;
  wire 140;
  wire 1400;
  wire 1401;
  wire 1402;
  wire 1403;
  wire 1404;
  wire 1405;
  wire 1406;
  wire 1407;
  wire 1408;
  wire 1409;
  wire 141;
  wire 1410;
  wire 1411;
  wire 1412;
  wire 1413;
  wire 1414;
  wire 1415;
  wire 1416;
  wire 1417;
  wire 1418;
  wire 1419;
  wire 142;
  wire 1420;
  wire 1421;
  wire 1422;
  wire 1423;
  wire 1424;
  wire 1425;
  wire 1426;
  wire 1427;
  wire 1428;
  wire 1429;
  wire 143;
  wire 1430;
  wire 1431;
  wire 1432;
  wire 1433;
  wire 1434;
  wire 1435;
  wire 1436;
  wire 1437;
  wire 1438;
  wire 1439;
  wire 144;
  wire 1440;
  wire 1441;
  wire 1442;
  wire 1443;
  wire 1444;
  wire 1445;
  wire 1446;
  wire 1447;
  wire 1448;
  wire 1449;
  wire 145;
  wire 1450;
  wire 1451;
  wire 1452;
  wire 1453;
  wire 1454;
  wire 1455;
  wire 1456;
  wire 1457;
  wire 1458;
  wire 1459;
  wire 146;
  wire 1460;
  wire 1461;
  wire 1462;
  wire 1463;
  wire 1464;
  wire 1465;
  wire 1466;
  wire 1467;
  wire 1468;
  wire 1469;
  wire 147;
  wire 1470;
  wire 1471;
  wire 1472;
  wire 1473;
  wire 1474;
  wire 1475;
  wire 1476;
  wire 1477;
  wire 1478;
  wire 1479;
  wire 148;
  wire 1480;
  wire 1481;
  wire 1482;
  wire 1483;
  wire 1484;
  wire 1485;
  wire 1486;
  wire 1487;
  wire 1488;
  wire 1489;
  wire 149;
  wire 1490;
  wire 1491;
  wire 1492;
  wire 1493;
  wire 1494;
  wire 1495;
  wire 1496;
  wire 1497;
  wire 1498;
  wire 1499;
  wire 150;
  wire 1500;
  wire 1501;
  wire 1502;
  wire 1503;
  wire 1504;
  wire 1505;
  wire 1506;
  wire 1507;
  wire 1508;
  wire 1509;
  wire 151;
  wire 1510;
  wire 1511;
  wire 1512;
  wire 1513;
  wire 1514;
  wire 1515;
  wire 1516;
  wire 1517;
  wire 1518;
  wire 1519;
  wire 152;
  wire 1520;
  wire 1521;
  wire 1522;
  wire 1523;
  wire 1524;
  wire 1525;
  wire 1526;
  wire 1527;
  wire 1528;
  wire 1529;
  wire 153;
  wire 1530;
  wire 1531;
  wire 1532;
  wire 1533;
  wire 1534;
  wire 1535;
  wire 1536;
  wire 1537;
  wire 1538;
  wire 1539;
  wire 154;
  wire 1540;
  wire 1541;
  wire 1542;
  wire 1543;
  wire 1544;
  wire 1545;
  wire 1546;
  wire 1547;
  wire 1548;
  wire 1549;
  wire 155;
  wire 1550;
  wire 1551;
  wire 1552;
  wire 1553;
  wire 1554;
  wire 1555;
  wire 1556;
  wire 1557;
  wire 1558;
  wire 1559;
  wire 156;
  wire 1560;
  wire 1561;
  wire 1562;
  wire 1563;
  wire 1564;
  wire 1565;
  wire 1566;
  wire 1567;
  wire 1568;
  wire 1569;
  wire 157;
  wire 1570;
  wire 1571;
  wire 1572;
  wire 1573;
  wire 1574;
  wire 1575;
  wire 1576;
  wire 1577;
  wire 1578;
  wire 1579;
  wire 158;
  wire 1580;
  wire 1581;
  wire 1582;
  wire 1583;
  wire 1584;
  wire 1585;
  wire 1586;
  wire 1587;
  wire 1588;
  wire 1589;
  wire 159;
  wire 1590;
  wire 1591;
  wire 1592;
  wire 1593;
  wire 1594;
  wire 1595;
  wire 1596;
  wire 1597;
  wire 1598;
  wire 1599;
  wire 160;
  wire 1600;
  wire 1601;
  wire 1602;
  wire 1603;
  wire 1604;
  wire 1605;
  wire 1606;
  wire 1607;
  wire 1608;
  wire 1609;
  wire 161;
  wire 1610;
  wire 1611;
  wire 1612;
  wire 1613;
  wire 1614;
  wire 1615;
  wire 1616;
  wire 1617;
  wire 1618;
  wire 1619;
  wire 162;
  wire 1620;
  wire 1621;
  wire 1622;
  wire 1623;
  wire 1624;
  wire 1625;
  wire 1626;
  wire 1627;
  wire 1628;
  wire 1629;
  wire 163;
  wire 1630;
  wire 1631;
  wire 1632;
  wire 1633;
  wire 1634;
  wire 1635;
  wire 1636;
  wire 1637;
  wire 1638;
  wire 1639;
  wire 164;
  wire 1640;
  wire 1641;
  wire 1642;
  wire 1643;
  wire 1644;
  wire 1645;
  wire 1646;
  wire 1647;
  wire 1648;
  wire 1649;
  wire 165;
  wire 1650;
  wire 1651;
  wire 1652;
  wire 1653;
  wire 1654;
  wire 1655;
  wire 1656;
  wire 1657;
  wire 1658;
  wire 1659;
  wire 166;
  wire 1660;
  wire 1661;
  wire 1662;
  wire 1663;
  wire 1664;
  wire 1665;
  wire 1666;
  wire 1667;
  wire 1668;
  wire 1669;
  wire 167;
  wire 1670;
  wire 1671;
  wire 1672;
  wire 1673;
  wire 1674;
  wire 1675;
  wire 1676;
  wire 1677;
  wire 1678;
  wire 1679;
  wire 168;
  wire 1680;
  wire 1681;
  wire 1682;
  wire 1683;
  wire 1684;
  wire 1685;
  wire 1686;
  wire 1687;
  wire 1688;
  wire 1689;
  wire 169;
  wire 1690;
  wire 1691;
  wire 1692;
  wire 1693;
  wire 1694;
  wire 1695;
  wire 1696;
  wire 1697;
  wire 1698;
  wire 1699;
  wire 170;
  wire 1700;
  wire 1701;
  wire 1702;
  wire 1703;
  wire 1704;
  wire 1705;
  wire 1706;
  wire 1707;
  wire 1708;
  wire 1709;
  wire 171;
  wire 1710;
  wire 1711;
  wire 1712;
  wire 1713;
  wire 1714;
  wire 1715;
  wire 1716;
  wire 1717;
  wire 1718;
  wire 1719;
  wire 172;
  wire 1720;
  wire 1721;
  wire 1722;
  wire 1723;
  wire 1724;
  wire 1725;
  wire 1726;
  wire 1727;
  wire 1728;
  wire 1729;
  wire 173;
  wire 1730;
  wire 1731;
  wire 1732;
  wire 1733;
  wire 1734;
  wire 1735;
  wire 1736;
  wire 1737;
  wire 1738;
  wire 1739;
  wire 174;
  wire 1740;
  wire 1741;
  wire 1742;
  wire 1743;
  wire 1744;
  wire 1745;
  wire 1746;
  wire 1747;
  wire 1748;
  wire 1749;
  wire 175;
  wire 1750;
  wire 1751;
  wire 1752;
  wire 1753;
  wire 1754;
  wire 1755;
  wire 1756;
  wire 1757;
  wire 1758;
  wire 1759;
  wire 176;
  wire 1760;
  wire 1761;
  wire 1762;
  wire 1763;
  wire 1764;
  wire 1765;
  wire 1766;
  wire 1767;
  wire 1768;
  wire 1769;
  wire 177;
  wire 1770;
  wire 1771;
  wire 1772;
  wire 1773;
  wire 1774;
  wire 1775;
  wire 1776;
  wire 1777;
  wire 1778;
  wire 1779;
  wire 178;
  wire 1780;
  wire 1781;
  wire 1782;
  wire 1783;
  wire 1784;
  wire 1785;
  wire 1786;
  wire 1787;
  wire 1788;
  wire 1789;
  wire 179;
  wire 1790;
  wire 1791;
  wire 1792;
  wire 1793;
  wire 1794;
  wire 1795;
  wire 1796;
  wire 1797;
  wire 1798;
  wire 1799;
  wire 180;
  wire 1800;
  wire 1801;
  wire 1802;
  wire 1803;
  wire 1804;
  wire 1805;
  wire 1806;
  wire 1807;
  wire 1808;
  wire 1809;
  wire 181;
  wire 1810;
  wire 1811;
  wire 1812;
  wire 1813;
  wire 1814;
  wire 1815;
  wire 1816;
  wire 1817;
  wire 1818;
  wire 1819;
  wire 182;
  wire 1820;
  wire 1821;
  wire 1822;
  wire 1823;
  wire 1824;
  wire 1825;
  wire 1826;
  wire 1827;
  wire 1828;
  wire 1829;
  wire 183;
  wire 1830;
  wire 1831;
  wire 1832;
  wire 1833;
  wire 1834;
  wire 1835;
  wire 1836;
  wire 1837;
  wire 1838;
  wire 1839;
  wire 184;
  wire 1840;
  wire 1841;
  wire 1842;
  wire 1843;
  wire 1844;
  wire 1845;
  wire 1846;
  wire 1847;
  wire 1848;
  wire 1849;
  wire 185;
  wire 1850;
  wire 1851;
  wire 1852;
  wire 1853;
  wire 1854;
  wire 1855;
  wire 1856;
  wire 1857;
  wire 1858;
  wire 1859;
  wire 186;
  wire 1860;
  wire 1861;
  wire 1862;
  wire 1863;
  wire 1864;
  wire 1865;
  wire 1866;
  wire 1867;
  wire 1868;
  wire 1869;
  wire 187;
  wire 1870;
  wire 1871;
  wire 1872;
  wire 1873;
  wire 1874;
  wire 1875;
  wire 1876;
  wire 1877;
  wire 1878;
  wire 1879;
  wire 188;
  wire 1880;
  wire 1881;
  wire 1882;
  wire 1883;
  wire 1884;
  wire 1885;
  wire 1886;
  wire 1887;
  wire 1888;
  wire 1889;
  wire 189;
  wire 1890;
  wire 1891;
  wire 1892;
  wire 1893;
  wire 1894;
  wire 1895;
  wire 1896;
  wire 1897;
  wire 1898;
  wire 1899;
  wire 190;
  wire 1900;
  wire 1901;
  wire 1902;
  wire 1903;
  wire 1904;
  wire 1905;
  wire 1906;
  wire 1907;
  wire 1908;
  wire 1909;
  wire 191;
  wire 1910;
  wire 1911;
  wire 1912;
  wire 1913;
  wire 1914;
  wire 1915;
  wire 1916;
  wire 1917;
  wire 1918;
  wire 1919;
  wire 192;
  wire 1920;
  wire 1921;
  wire 1922;
  wire 1923;
  wire 1924;
  wire 1925;
  wire 1926;
  wire 1927;
  wire 1928;
  wire 1929;
  wire 193;
  wire 1930;
  wire 1931;
  wire 1932;
  wire 1933;
  wire 1934;
  wire 1935;
  wire 1936;
  wire 1937;
  wire 1938;
  wire 1939;
  wire 194;
  wire 1940;
  wire 1941;
  wire 1942;
  wire 1943;
  wire 1944;
  wire 1945;
  wire 1946;
  wire 1947;
  wire 1948;
  wire 1949;
  wire 195;
  wire 1950;
  wire 1951;
  wire 1952;
  wire 1953;
  wire 1954;
  wire 1955;
  wire 1956;
  wire 1957;
  wire 1958;
  wire 1959;
  wire 196;
  wire 1960;
  wire 1961;
  wire 1962;
  wire 1963;
  wire 1964;
  wire 1965;
  wire 1966;
  wire 1967;
  wire 1968;
  wire 1969;
  wire 197;
  wire 1970;
  wire 1971;
  wire 1972;
  wire 1973;
  wire 1974;
  wire 1975;
  wire 1976;
  wire 1977;
  wire 1978;
  wire 1979;
  wire 198;
  wire 1980;
  wire 1981;
  wire 1982;
  wire 1983;
  wire 1984;
  wire 1985;
  wire 1986;
  wire 1987;
  wire 1988;
  wire 1989;
  wire 199;
  wire 1990;
  wire 1991;
  wire 1992;
  wire 1993;
  wire 1994;
  wire 1995;
  wire 1996;
  wire 1997;
  wire 1998;
  wire 1999;
  wire 2;
  wire 20;
  wire 200;
  wire 2000;
  wire 2001;
  wire 2002;
  wire 2003;
  wire 2004;
  wire 2005;
  wire 2006;
  wire 2007;
  wire 2008;
  wire 2009;
  wire 201;
  wire 2010;
  wire 2011;
  wire 2012;
  wire 2013;
  wire 2014;
  wire 2015;
  wire 2016;
  wire 2017;
  wire 2018;
  wire 2019;
  wire 202;
  wire 2020;
  wire 2021;
  wire 2022;
  wire 2023;
  wire 2024;
  wire 2025;
  wire 2026;
  wire 2027;
  wire 2028;
  wire 2029;
  wire 203;
  wire 2030;
  wire 2031;
  wire 2032;
  wire 2033;
  wire 2034;
  wire 2035;
  wire 2036;
  wire 2037;
  wire 2038;
  wire 2039;
  wire 204;
  wire 2040;
  wire 2041;
  wire 2042;
  wire 2043;
  wire 2044;
  wire 2045;
  wire 2046;
  wire 2047;
  wire 2048;
  wire 2049;
  wire 205;
  wire 2050;
  wire 2051;
  wire 2052;
  wire 2053;
  wire 2054;
  wire 2055;
  wire 2056;
  wire 2057;
  wire 2058;
  wire 2059;
  wire 206;
  wire 2060;
  wire 2061;
  wire 2062;
  wire 2063;
  wire 2064;
  wire 2065;
  wire 2066;
  wire 2067;
  wire 2068;
  wire 2069;
  wire 207;
  wire 2070;
  wire 2071;
  wire 2072;
  wire 2073;
  wire 2074;
  wire 2075;
  wire 2076;
  wire 2077;
  wire 2078;
  wire 2079;
  wire 208;
  wire 2080;
  wire 2081;
  wire 2082;
  wire 2083;
  wire 2084;
  wire 2085;
  wire 2086;
  wire 2087;
  wire 2088;
  wire 2089;
  wire 209;
  wire 2090;
  wire 2091;
  wire 2092;
  wire 2093;
  wire 2094;
  wire 2095;
  wire 2096;
  wire 2097;
  wire 2098;
  wire 2099;
  wire 21;
  wire 210;
  wire 2100;
  wire 2101;
  wire 2102;
  wire 2103;
  wire 2104;
  wire 2105;
  wire 2106;
  wire 2107;
  wire 2108;
  wire 2109;
  wire 211;
  wire 2110;
  wire 2111;
  wire 2112;
  wire 2113;
  wire 2114;
  wire 2115;
  wire 2116;
  wire 2117;
  wire 2118;
  wire 2119;
  wire 212;
  wire 2120;
  wire 2121;
  wire 2122;
  wire 2123;
  wire 2124;
  wire 2125;
  wire 2126;
  wire 2127;
  wire 2128;
  wire 2129;
  wire 213;
  wire 2130;
  wire 2131;
  wire 2132;
  wire 2133;
  wire 2134;
  wire 2135;
  wire 2136;
  wire 2137;
  wire 2138;
  wire 2139;
  wire 214;
  wire 2140;
  wire 2141;
  wire 2142;
  wire 2143;
  wire 2144;
  wire 2145;
  wire 2146;
  wire 2147;
  wire 2148;
  wire 2149;
  wire 215;
  wire 2150;
  wire 2151;
  wire 2152;
  wire 2153;
  wire 2154;
  wire 2155;
  wire 2156;
  wire 2157;
  wire 2158;
  wire 2159;
  wire 216;
  wire 2160;
  wire 2161;
  wire 2162;
  wire 2163;
  wire 2164;
  wire 2165;
  wire 2166;
  wire 2167;
  wire 2168;
  wire 2169;
  wire 217;
  wire 2170;
  wire 2171;
  wire 2172;
  wire 2173;
  wire 2174;
  wire 2175;
  wire 2176;
  wire 2177;
  wire 2178;
  wire 2179;
  wire 218;
  wire 2180;
  wire 2181;
  wire 2182;
  wire 2183;
  wire 2184;
  wire 2185;
  wire 2186;
  wire 2187;
  wire 2188;
  wire 2189;
  wire 219;
  wire 2190;
  wire 2191;
  wire 2192;
  wire 2193;
  wire 2194;
  wire 2195;
  wire 2196;
  wire 2197;
  wire 2198;
  wire 2199;
  wire 22;
  wire 220;
  wire 2200;
  wire 2201;
  wire 2202;
  wire 2203;
  wire 2204;
  wire 2205;
  wire 2206;
  wire 2207;
  wire 2208;
  wire 2209;
  wire 221;
  wire 2210;
  wire 2211;
  wire 2212;
  wire 2213;
  wire 2214;
  wire 2215;
  wire 2216;
  wire 2217;
  wire 2218;
  wire 2219;
  wire 222;
  wire 2220;
  wire 2221;
  wire 2222;
  wire 2223;
  wire 2224;
  wire 2225;
  wire 2226;
  wire 2227;
  wire 2228;
  wire 2229;
  wire 223;
  wire 2230;
  wire 2231;
  wire 2232;
  wire 2233;
  wire 2234;
  wire 2235;
  wire 2236;
  wire 2237;
  wire 2238;
  wire 2239;
  wire 224;
  wire 2240;
  wire 2241;
  wire 2242;
  wire 2243;
  wire 2244;
  wire 2245;
  wire 2246;
  wire 2247;
  wire 2248;
  wire 2249;
  wire 225;
  wire 2250;
  wire 2251;
  wire 2252;
  wire 2253;
  wire 2254;
  wire 2255;
  wire 2256;
  wire 2257;
  wire 2258;
  wire 2259;
  wire 226;
  wire 2260;
  wire 2261;
  wire 2262;
  wire 2263;
  wire 2264;
  wire 2265;
  wire 2266;
  wire 2267;
  wire 2268;
  wire 2269;
  wire 227;
  wire 2270;
  wire 2271;
  wire 2272;
  wire 2273;
  wire 2274;
  wire 2275;
  wire 2276;
  wire 2277;
  wire 2278;
  wire 2279;
  wire 228;
  wire 2280;
  wire 2281;
  wire 2282;
  wire 2283;
  wire 2284;
  wire 2285;
  wire 2286;
  wire 2287;
  wire 2288;
  wire 2289;
  wire 229;
  wire 2290;
  wire 2291;
  wire 2292;
  wire 2293;
  wire 2294;
  wire 2295;
  wire 2296;
  wire 2297;
  wire 2298;
  wire 2299;
  wire 23;
  wire 230;
  wire 2300;
  wire 2301;
  wire 2302;
  wire 2303;
  wire 2304;
  wire 2305;
  wire 2306;
  wire 2307;
  wire 2308;
  wire 2309;
  wire 231;
  wire 2310;
  wire 2311;
  wire 2312;
  wire 2313;
  wire 2314;
  wire 2315;
  wire 2316;
  wire 2317;
  wire 2318;
  wire 2319;
  wire 232;
  wire 2320;
  wire 2321;
  wire 2322;
  wire 2323;
  wire 2324;
  wire 2325;
  wire 2326;
  wire 2327;
  wire 2328;
  wire 2329;
  wire 233;
  wire 2330;
  wire 2331;
  wire 2332;
  wire 2333;
  wire 2334;
  wire 2335;
  wire 2336;
  wire 2337;
  wire 2338;
  wire 2339;
  wire 234;
  wire 2340;
  wire 2341;
  wire 2342;
  wire 2343;
  wire 2344;
  wire 2345;
  wire 2346;
  wire 2347;
  wire 2348;
  wire 2349;
  wire 235;
  wire 2350;
  wire 2351;
  wire 2352;
  wire 2353;
  wire 2354;
  wire 2355;
  wire 2356;
  wire 2357;
  wire 2358;
  wire 2359;
  wire 236;
  wire 2360;
  wire 2361;
  wire 2362;
  wire 2363;
  wire 2364;
  wire 2365;
  wire 2366;
  wire 2367;
  wire 2368;
  wire 2369;
  wire 237;
  wire 2370;
  wire 2371;
  wire 2372;
  wire 2373;
  wire 2374;
  wire 2375;
  wire 2376;
  wire 2377;
  wire 2378;
  wire 2379;
  wire 238;
  wire 2380;
  wire 2381;
  wire 2382;
  wire 2383;
  wire 2384;
  wire 2385;
  wire 2386;
  wire 2387;
  wire 2388;
  wire 2389;
  wire 239;
  wire 2390;
  wire 2391;
  wire 2392;
  wire 2393;
  wire 2394;
  wire 2395;
  wire 2396;
  wire 2397;
  wire 2398;
  wire 2399;
  wire 24;
  wire 240;
  wire 2400;
  wire 2401;
  wire 2402;
  wire 2403;
  wire 2404;
  wire 2405;
  wire 2406;
  wire 2407;
  wire 2408;
  wire 2409;
  wire 241;
  wire 2410;
  wire 2411;
  wire 2412;
  wire 2413;
  wire 2414;
  wire 2415;
  wire 2416;
  wire 2417;
  wire 2418;
  wire 2419;
  wire 242;
  wire 2420;
  wire 2421;
  wire 2422;
  wire 2423;
  wire 2424;
  wire 2425;
  wire 2426;
  wire 2427;
  wire 2428;
  wire 2429;
  wire 243;
  wire 2430;
  wire 2431;
  wire 2432;
  wire 2433;
  wire 2434;
  wire 2435;
  wire 2436;
  wire 2437;
  wire 2438;
  wire 2439;
  wire 244;
  wire 2440;
  wire 2441;
  wire 2442;
  wire 2443;
  wire 2444;
  wire 2445;
  wire 2446;
  wire 2447;
  wire 2448;
  wire 2449;
  wire 245;
  wire 2450;
  wire 2451;
  wire 2452;
  wire 2453;
  wire 2454;
  wire 2455;
  wire 2456;
  wire 2457;
  wire 2458;
  wire 2459;
  wire 246;
  wire 2460;
  wire 2461;
  wire 2462;
  wire 2463;
  wire 2464;
  wire 2465;
  wire 2466;
  wire 2467;
  wire 2468;
  wire 2469;
  wire 247;
  wire 2470;
  wire 2471;
  wire 2472;
  wire 2473;
  wire 2474;
  wire 2475;
  wire 2476;
  wire 2477;
  wire 2478;
  wire 2479;
  wire 248;
  wire 2480;
  wire 2481;
  wire 2482;
  wire 2483;
  wire 2484;
  wire 2485;
  wire 2486;
  wire 2487;
  wire 2488;
  wire 2489;
  wire 249;
  wire 2490;
  wire 2491;
  wire 2492;
  wire 2493;
  wire 2494;
  wire 2495;
  wire 2496;
  wire 2497;
  wire 2498;
  wire 2499;
  wire 25;
  wire 250;
  wire 2500;
  wire 2501;
  wire 2502;
  wire 2503;
  wire 2504;
  wire 2505;
  wire 2506;
  wire 2507;
  wire 2508;
  wire 2509;
  wire 251;
  wire 2510;
  wire 2511;
  wire 2512;
  wire 2513;
  wire 2514;
  wire 2515;
  wire 2516;
  wire 2517;
  wire 2518;
  wire 2519;
  wire 252;
  wire 2520;
  wire 2521;
  wire 2522;
  wire 2523;
  wire 2524;
  wire 2525;
  wire 2526;
  wire 2527;
  wire 2528;
  wire 2529;
  wire 253;
  wire 2530;
  wire 2531;
  wire 2532;
  wire 2533;
  wire 2534;
  wire 2535;
  wire 2536;
  wire 2537;
  wire 2538;
  wire 2539;
  wire 254;
  wire 2540;
  wire 2541;
  wire 2542;
  wire 2543;
  wire 2544;
  wire 2545;
  wire 2546;
  wire 2547;
  wire 2548;
  wire 2549;
  wire 255;
  wire 2550;
  wire 2551;
  wire 2552;
  wire 2553;
  wire 2554;
  wire 2555;
  wire 2556;
  wire 2557;
  wire 2558;
  wire 2559;
  wire 256;
  wire 2560;
  wire 2561;
  wire 2562;
  wire 2563;
  wire 2564;
  wire 2565;
  wire 2566;
  wire 2567;
  wire 2568;
  wire 2569;
  wire 257;
  wire 2570;
  wire 2571;
  wire 2572;
  wire 2573;
  wire 2574;
  wire 2575;
  wire 2576;
  wire 2577;
  wire 2578;
  wire 2579;
  wire 258;
  wire 2580;
  wire 2581;
  wire 2582;
  wire 2583;
  wire 2584;
  wire 2585;
  wire 2586;
  wire 2587;
  wire 2588;
  wire 2589;
  wire 259;
  wire 2590;
  wire 2591;
  wire 2592;
  wire 2593;
  wire 2594;
  wire 2595;
  wire 2596;
  wire 2597;
  wire 2598;
  wire 2599;
  wire 26;
  wire 260;
  wire 2600;
  wire 2601;
  wire 2602;
  wire 2603;
  wire 2604;
  wire 2605;
  wire 2606;
  wire 2607;
  wire 2608;
  wire 2609;
  wire 261;
  wire 2610;
  wire 2611;
  wire 2612;
  wire 2613;
  wire 2614;
  wire 2615;
  wire 2616;
  wire 2617;
  wire 2618;
  wire 2619;
  wire 262;
  wire 2620;
  wire 2621;
  wire 2622;
  wire 2623;
  wire 2624;
  wire 2625;
  wire 2626;
  wire 2627;
  wire 2628;
  wire 2629;
  wire 263;
  wire 2630;
  wire 2631;
  wire 2632;
  wire 2633;
  wire 2634;
  wire 2635;
  wire 2636;
  wire 2637;
  wire 2638;
  wire 2639;
  wire 264;
  wire 2640;
  wire 2641;
  wire 2642;
  wire 2643;
  wire 2644;
  wire 2645;
  wire 2646;
  wire 2647;
  wire 2648;
  wire 2649;
  wire 265;
  wire 2650;
  wire 2651;
  wire 2652;
  wire 2653;
  wire 2654;
  wire 2655;
  wire 2656;
  wire 2657;
  wire 2658;
  wire 2659;
  wire 266;
  wire 2660;
  wire 2661;
  wire 2662;
  wire 2663;
  wire 2664;
  wire 2665;
  wire 2666;
  wire 2667;
  wire 2668;
  wire 2669;
  wire 267;
  wire 2670;
  wire 2671;
  wire 2672;
  wire 2673;
  wire 2674;
  wire 2675;
  wire 2676;
  wire 2677;
  wire 2678;
  wire 2679;
  wire 268;
  wire 2680;
  wire 2681;
  wire 2682;
  wire 2683;
  wire 2684;
  wire 2685;
  wire 2686;
  wire 2687;
  wire 2688;
  wire 2689;
  wire 269;
  wire 2690;
  wire 2691;
  wire 2692;
  wire 2693;
  wire 2694;
  wire 2695;
  wire 2696;
  wire 2697;
  wire 2698;
  wire 2699;
  wire 27;
  wire 270;
  wire 2700;
  wire 2701;
  wire 2702;
  wire 2703;
  wire 2704;
  wire 2705;
  wire 2706;
  wire 2707;
  wire 2708;
  wire 2709;
  wire 271;
  wire 2710;
  wire 2711;
  wire 2712;
  wire 2713;
  wire 2714;
  wire 2715;
  wire 2716;
  wire 2717;
  wire 2718;
  wire 2719;
  wire 272;
  wire 2720;
  wire 2721;
  wire 2722;
  wire 2723;
  wire 2724;
  wire 2725;
  wire 2726;
  wire 2727;
  wire 2728;
  wire 2729;
  wire 273;
  wire 2730;
  wire 2731;
  wire 2732;
  wire 2733;
  wire 2734;
  wire 2735;
  wire 2736;
  wire 2737;
  wire 2738;
  wire 2739;
  wire 274;
  wire 2740;
  wire 2741;
  wire 2742;
  wire 2743;
  wire 2744;
  wire 2745;
  wire 2746;
  wire 2747;
  wire 2748;
  wire 2749;
  wire 275;
  wire 2750;
  wire 2751;
  wire 2752;
  wire 2753;
  wire 2754;
  wire 2755;
  wire 2756;
  wire 2757;
  wire 2758;
  wire 2759;
  wire 276;
  wire 2760;
  wire 2761;
  wire 2762;
  wire 2763;
  wire 2764;
  wire 2765;
  wire 2766;
  wire 2767;
  wire 2768;
  wire 2769;
  wire 277;
  wire 2770;
  wire 2771;
  wire 2772;
  wire 2773;
  wire 2774;
  wire 2775;
  wire 2776;
  wire 2777;
  wire 2778;
  wire 2779;
  wire 278;
  wire 2780;
  wire 2781;
  wire 2782;
  wire 2783;
  wire 2784;
  wire 2785;
  wire 2786;
  wire 2787;
  wire 2788;
  wire 2789;
  wire 279;
  wire 2790;
  wire 2791;
  wire 2792;
  wire 2793;
  wire 2794;
  wire 2795;
  wire 2796;
  wire 2797;
  wire 2798;
  wire 2799;
  wire 280;
  wire 2800;
  wire 2801;
  wire 2802;
  wire 2803;
  wire 2804;
  wire 2805;
  wire 2806;
  wire 2807;
  wire 2808;
  wire 2809;
  wire 281;
  wire 2810;
  wire 2811;
  wire 2812;
  wire 2813;
  wire 2814;
  wire 2815;
  wire 2816;
  wire 2817;
  wire 2818;
  wire 2819;
  wire 282;
  wire 2820;
  wire 2821;
  wire 2822;
  wire 2823;
  wire 2824;
  wire 2825;
  wire 2826;
  wire 2827;
  wire 2828;
  wire 2829;
  wire 283;
  wire 2830;
  wire 2831;
  wire 2832;
  wire 2833;
  wire 2834;
  wire 2835;
  wire 2836;
  wire 2837;
  wire 2838;
  wire 2839;
  wire 284;
  wire 2840;
  wire 2841;
  wire 2842;
  wire 2843;
  wire 2844;
  wire 2845;
  wire 2846;
  wire 2847;
  wire 2848;
  wire 2849;
  wire 285;
  wire 2850;
  wire 2851;
  wire 2852;
  wire 2853;
  wire 2854;
  wire 2855;
  wire 2856;
  wire 2857;
  wire 2858;
  wire 2859;
  wire 286;
  wire 2860;
  wire 2861;
  wire 2862;
  wire 2863;
  wire 2864;
  wire 2865;
  wire 2866;
  wire 2867;
  wire 2868;
  wire 2869;
  wire 287;
  wire 2870;
  wire 2871;
  wire 2872;
  wire 2873;
  wire 2874;
  wire 2875;
  wire 2876;
  wire 2877;
  wire 2878;
  wire 2879;
  wire 288;
  wire 2880;
  wire 2881;
  wire 2882;
  wire 2883;
  wire 2884;
  wire 2885;
  wire 2886;
  wire 2887;
  wire 2888;
  wire 2889;
  wire 289;
  wire 2890;
  wire 2891;
  wire 2892;
  wire 2893;
  wire 2894;
  wire 2895;
  wire 2896;
  wire 2897;
  wire 2898;
  wire 2899;
  wire 290;
  wire 2900;
  wire 2901;
  wire 2902;
  wire 2903;
  wire 2904;
  wire 2905;
  wire 2906;
  wire 2907;
  wire 2908;
  wire 2909;
  wire 291;
  wire 2910;
  wire 2911;
  wire 2912;
  wire 2913;
  wire 2914;
  wire 2915;
  wire 2916;
  wire 2917;
  wire 2918;
  wire 2919;
  wire 292;
  wire 2920;
  wire 2921;
  wire 2922;
  wire 2923;
  wire 2924;
  wire 2925;
  wire 2926;
  wire 2927;
  wire 2928;
  wire 2929;
  wire 293;
  wire 2930;
  wire 2931;
  wire 2932;
  wire 2933;
  wire 2934;
  wire 2935;
  wire 2936;
  wire 2937;
  wire 2938;
  wire 2939;
  wire 294;
  wire 2940;
  wire 2941;
  wire 2942;
  wire 2943;
  wire 2944;
  wire 2945;
  wire 2946;
  wire 2947;
  wire 2948;
  wire 2949;
  wire 295;
  wire 2950;
  wire 2951;
  wire 2952;
  wire 2953;
  wire 2954;
  wire 2955;
  wire 2956;
  wire 2957;
  wire 2958;
  wire 2959;
  wire 296;
  wire 2960;
  wire 2961;
  wire 2962;
  wire 2963;
  wire 2964;
  wire 2965;
  wire 2966;
  wire 2967;
  wire 2968;
  wire 2969;
  wire 297;
  wire 2970;
  wire 2971;
  wire 2972;
  wire 2973;
  wire 2974;
  wire 2975;
  wire 2976;
  wire 2977;
  wire 2978;
  wire 2979;
  wire 298;
  wire 2980;
  wire 2981;
  wire 2982;
  wire 2983;
  wire 2984;
  wire 2985;
  wire 2986;
  wire 2987;
  wire 2988;
  wire 2989;
  wire 299;
  wire 2990;
  wire 2991;
  wire 2992;
  wire 2993;
  wire 2994;
  wire 2995;
  wire 2996;
  wire 2997;
  wire 2998;
  wire 2999;
  wire 3;
  wire 300;
  wire 3000;
  wire 3001;
  wire 3002;
  wire 3003;
  wire 3004;
  wire 3005;
  wire 3006;
  wire 3007;
  wire 3008;
  wire 3009;
  wire 301;
  wire 3010;
  wire 3011;
  wire 3012;
  wire 3013;
  wire 3014;
  wire 3015;
  wire 3016;
  wire 3017;
  wire 3018;
  wire 3019;
  wire 302;
  wire 3020;
  wire 3021;
  wire 3022;
  wire 3023;
  wire 3024;
  wire 3025;
  wire 3026;
  wire 3027;
  wire 3028;
  wire 3029;
  wire 303;
  wire 3030;
  wire 3031;
  wire 3032;
  wire 3033;
  wire 3034;
  wire 3035;
  wire 3036;
  wire 3037;
  wire 3038;
  wire 3039;
  wire 304;
  wire 3040;
  wire 3041;
  wire 3042;
  wire 3043;
  wire 3044;
  wire 3045;
  wire 3046;
  wire 3047;
  wire 3048;
  wire 3049;
  wire 305;
  wire 3050;
  wire 3051;
  wire 3052;
  wire 3053;
  wire 3054;
  wire 3055;
  wire 3056;
  wire 3057;
  wire 3058;
  wire 3059;
  wire 306;
  wire 3060;
  wire 3061;
  wire 3062;
  wire 3063;
  wire 3064;
  wire 3065;
  wire 3066;
  wire 3067;
  wire 3068;
  wire 3069;
  wire 307;
  wire 3070;
  wire 3071;
  wire 3072;
  wire 3073;
  wire 3074;
  wire 3075;
  wire 3076;
  wire 3077;
  wire 3078;
  wire 3079;
  wire 308;
  wire 3080;
  wire 3081;
  wire 3082;
  wire 3083;
  wire 3084;
  wire 3085;
  wire 3086;
  wire 3087;
  wire 309;
  wire 310;
  wire 311;
  wire 312;
  wire 313;
  wire 314;
  wire 315;
  wire 316;
  wire 317;
  wire 318;
  wire 319;
  wire 320;
  wire 321;
  wire 322;
  wire 323;
  wire 324;
  wire 325;
  wire 326;
  wire 327;
  wire 328;
  wire 329;
  wire 330;
  wire 331;
  wire 332;
  wire 333;
  wire 334;
  wire 335;
  wire 336;
  wire 337;
  wire 338;
  wire 339;
  wire 340;
  wire 341;
  wire 342;
  wire 343;
  wire 344;
  wire 345;
  wire 346;
  wire 347;
  wire 348;
  wire 349;
  wire 350;
  wire 351;
  wire 352;
  wire 353;
  wire 354;
  wire 355;
  wire 356;
  wire 357;
  wire 358;
  wire 359;
  wire 360;
  wire 361;
  wire 362;
  wire 363;
  wire 364;
  wire 365;
  wire 366;
  wire 367;
  wire 368;
  wire 369;
  wire 37;
  wire 370;
  wire 371;
  wire 372;
  wire 373;
  wire 374;
  wire 375;
  wire 376;
  wire 377;
  wire 378;
  wire 379;
  wire 38;
  wire 380;
  wire 381;
  wire 382;
  wire 383;
  wire 384;
  wire 385;
  wire 386;
  wire 387;
  wire 388;
  wire 389;
  wire 39;
  wire 390;
  wire 391;
  wire 392;
  wire 393;
  wire 394;
  wire 395;
  wire 396;
  wire 397;
  wire 398;
  wire 399;
  wire 400;
  wire 401;
  wire 402;
  wire 403;
  wire 404;
  wire 405;
  wire 406;
  wire 407;
  wire 408;
  wire 409;
  wire 410;
  wire 411;
  wire 412;
  wire 413;
  wire 414;
  wire 415;
  wire 416;
  wire 417;
  wire 418;
  wire 419;
  wire 420;
  wire 421;
  wire 422;
  wire 423;
  wire 424;
  wire 425;
  wire 426;
  wire 427;
  wire 428;
  wire 429;
  wire 430;
  wire 431;
  wire 432;
  wire 433;
  wire 434;
  wire 435;
  wire 436;
  wire 437;
  wire 438;
  wire 439;
  wire 44;
  wire 440;
  wire 441;
  wire 442;
  wire 443;
  wire 444;
  wire 445;
  wire 446;
  wire 447;
  wire 448;
  wire 449;
  wire 45;
  wire 450;
  wire 451;
  wire 452;
  wire 453;
  wire 454;
  wire 455;
  wire 456;
  wire 457;
  wire 458;
  wire 459;
  wire 46;
  wire 460;
  wire 461;
  wire 462;
  wire 463;
  wire 464;
  wire 465;
  wire 466;
  wire 467;
  wire 468;
  wire 469;
  wire 47;
  wire 470;
  wire 471;
  wire 472;
  wire 473;
  wire 474;
  wire 475;
  wire 476;
  wire 477;
  wire 478;
  wire 479;
  wire 48;
  wire 480;
  wire 481;
  wire 482;
  wire 483;
  wire 484;
  wire 485;
  wire 486;
  wire 487;
  wire 488;
  wire 489;
  wire 49;
  wire 490;
  wire 491;
  wire 492;
  wire 493;
  wire 494;
  wire 495;
  wire 496;
  wire 497;
  wire 498;
  wire 499;
  wire 50;
  wire 500;
  wire 501;
  wire 502;
  wire 503;
  wire 504;
  wire 505;
  wire 506;
  wire 507;
  wire 508;
  wire 509;
  wire 51;
  wire 510;
  wire 511;
  wire 512;
  wire 513;
  wire 514;
  wire 515;
  wire 516;
  wire 517;
  wire 518;
  wire 519;
  wire 52;
  wire 520;
  wire 521;
  wire 522;
  wire 523;
  wire 524;
  wire 525;
  wire 526;
  wire 527;
  wire 528;
  wire 529;
  wire 53;
  wire 530;
  wire 531;
  wire 532;
  wire 533;
  wire 534;
  wire 535;
  wire 536;
  wire 537;
  wire 538;
  wire 539;
  wire 54;
  wire 540;
  wire 541;
  wire 542;
  wire 543;
  wire 544;
  wire 545;
  wire 546;
  wire 547;
  wire 548;
  wire 549;
  wire 55;
  wire 550;
  wire 551;
  wire 552;
  wire 553;
  wire 554;
  wire 555;
  wire 556;
  wire 557;
  wire 558;
  wire 559;
  wire 56;
  wire 560;
  wire 561;
  wire 562;
  wire 563;
  wire 564;
  wire 565;
  wire 566;
  wire 567;
  wire 568;
  wire 569;
  wire 57;
  wire 570;
  wire 571;
  wire 572;
  wire 573;
  wire 574;
  wire 575;
  wire 576;
  wire 577;
  wire 578;
  wire 579;
  wire 58;
  wire 580;
  wire 581;
  wire 582;
  wire 583;
  wire 584;
  wire 585;
  wire 586;
  wire 587;
  wire 588;
  wire 589;
  wire 59;
  wire 590;
  wire 591;
  wire 592;
  wire 593;
  wire 594;
  wire 595;
  wire 596;
  wire 597;
  wire 598;
  wire 599;
  wire 60;
  wire 600;
  wire 601;
  wire 602;
  wire 603;
  wire 604;
  wire 605;
  wire 606;
  wire 607;
  wire 608;
  wire 609;
  wire 61;
  wire 610;
  wire 611;
  wire 612;
  wire 613;
  wire 614;
  wire 615;
  wire 616;
  wire 617;
  wire 618;
  wire 619;
  wire 62;
  wire 620;
  wire 621;
  wire 622;
  wire 623;
  wire 624;
  wire 625;
  wire 626;
  wire 627;
  wire 628;
  wire 629;
  wire 63;
  wire 630;
  wire 631;
  wire 632;
  wire 633;
  wire 634;
  wire 635;
  wire 636;
  wire 637;
  wire 638;
  wire 639;
  wire 64;
  wire 640;
  wire 641;
  wire 642;
  wire 643;
  wire 644;
  wire 645;
  wire 646;
  wire 647;
  wire 648;
  wire 649;
  wire 65;
  wire 650;
  wire 651;
  wire 652;
  wire 653;
  wire 654;
  wire 655;
  wire 656;
  wire 657;
  wire 658;
  wire 659;
  wire 66;
  wire 660;
  wire 661;
  wire 662;
  wire 663;
  wire 664;
  wire 665;
  wire 666;
  wire 667;
  wire 668;
  wire 669;
  wire 67;
  wire 670;
  wire 671;
  wire 672;
  wire 673;
  wire 674;
  wire 675;
  wire 676;
  wire 677;
  wire 678;
  wire 679;
  wire 68;
  wire 680;
  wire 681;
  wire 682;
  wire 683;
  wire 684;
  wire 685;
  wire 686;
  wire 687;
  wire 688;
  wire 689;
  wire 69;
  wire 690;
  wire 691;
  wire 692;
  wire 693;
  wire 694;
  wire 695;
  wire 696;
  wire 697;
  wire 698;
  wire 699;
  wire 70;
  wire 700;
  wire 701;
  wire 702;
  wire 703;
  wire 704;
  wire 705;
  wire 706;
  wire 707;
  wire 708;
  wire 709;
  wire 71;
  wire 710;
  wire 711;
  wire 712;
  wire 713;
  wire 714;
  wire 715;
  wire 716;
  wire 717;
  wire 718;
  wire 719;
  wire 72;
  wire 720;
  wire 721;
  wire 722;
  wire 723;
  wire 724;
  wire 725;
  wire 726;
  wire 727;
  wire 728;
  wire 729;
  wire 73;
  wire 730;
  wire 731;
  wire 732;
  wire 733;
  wire 734;
  wire 735;
  wire 736;
  wire 737;
  wire 738;
  wire 739;
  wire 74;
  wire 740;
  wire 741;
  wire 742;
  wire 743;
  wire 744;
  wire 745;
  wire 746;
  wire 747;
  wire 748;
  wire 749;
  wire 75;
  wire 750;
  wire 751;
  wire 752;
  wire 753;
  wire 754;
  wire 755;
  wire 756;
  wire 757;
  wire 758;
  wire 759;
  wire 76;
  wire 760;
  wire 761;
  wire 762;
  wire 763;
  wire 764;
  wire 765;
  wire 766;
  wire 767;
  wire 768;
  wire 769;
  wire 77;
  wire 770;
  wire 771;
  wire 772;
  wire 773;
  wire 774;
  wire 775;
  wire 776;
  wire 777;
  wire 778;
  wire 779;
  wire 78;
  wire 780;
  wire 781;
  wire 782;
  wire 783;
  wire 784;
  wire 785;
  wire 786;
  wire 787;
  wire 788;
  wire 789;
  wire 79;
  wire 790;
  wire 791;
  wire 792;
  wire 793;
  wire 794;
  wire 795;
  wire 796;
  wire 797;
  wire 798;
  wire 799;
  wire 80;
  wire 800;
  wire 801;
  wire 802;
  wire 803;
  wire 804;
  wire 805;
  wire 806;
  wire 807;
  wire 808;
  wire 809;
  wire 81;
  wire 810;
  wire 811;
  wire 812;
  wire 813;
  wire 814;
  wire 815;
  wire 816;
  wire 817;
  wire 818;
  wire 819;
  wire 82;
  wire 820;
  wire 821;
  wire 822;
  wire 823;
  wire 824;
  wire 825;
  wire 826;
  wire 827;
  wire 828;
  wire 829;
  wire 83;
  wire 830;
  wire 831;
  wire 832;
  wire 833;
  wire 834;
  wire 835;
  wire 836;
  wire 837;
  wire 838;
  wire 839;
  wire 84;
  wire 840;
  wire 841;
  wire 842;
  wire 843;
  wire 844;
  wire 845;
  wire 846;
  wire 847;
  wire 848;
  wire 849;
  wire 85;
  wire 850;
  wire 851;
  wire 852;
  wire 853;
  wire 854;
  wire 855;
  wire 856;
  wire 857;
  wire 858;
  wire 859;
  wire 86;
  wire 860;
  wire 861;
  wire 862;
  wire 863;
  wire 864;
  wire 865;
  wire 866;
  wire 867;
  wire 868;
  wire 869;
  wire 87;
  wire 870;
  wire 871;
  wire 872;
  wire 873;
  wire 874;
  wire 875;
  wire 876;
  wire 877;
  wire 878;
  wire 879;
  wire 88;
  wire 880;
  wire 881;
  wire 882;
  wire 883;
  wire 884;
  wire 885;
  wire 886;
  wire 887;
  wire 888;
  wire 889;
  wire 89;
  wire 890;
  wire 891;
  wire 892;
  wire 893;
  wire 894;
  wire 895;
  wire 896;
  wire 897;
  wire 898;
  wire 899;
  wire 90;
  wire 900;
  wire 901;
  wire 902;
  wire 903;
  wire 904;
  wire 905;
  wire 906;
  wire 907;
  wire 908;
  wire 909;
  wire 91;
  wire 910;
  wire 911;
  wire 912;
  wire 913;
  wire 914;
  wire 915;
  wire 916;
  wire 917;
  wire 918;
  wire 919;
  wire 92;
  wire 920;
  wire 921;
  wire 922;
  wire 923;
  wire 924;
  wire 925;
  wire 926;
  wire 927;
  wire 928;
  wire 929;
  wire 93;
  wire 930;
  wire 931;
  wire 932;
  wire 933;
  wire 934;
  wire 935;
  wire 936;
  wire 937;
  wire 938;
  wire 939;
  wire 94;
  wire 940;
  wire 941;
  wire 942;
  wire 943;
  wire 944;
  wire 945;
  wire 946;
  wire 947;
  wire 948;
  wire 949;
  wire 95;
  wire 950;
  wire 951;
  wire 952;
  wire 953;
  wire 954;
  wire 955;
  wire 956;
  wire 957;
  wire 958;
  wire 959;
  wire 96;
  wire 960;
  wire 961;
  wire 962;
  wire 963;
  wire 964;
  wire 965;
  wire 966;
  wire 967;
  wire 968;
  wire 969;
  wire 97;
  wire 970;
  wire 971;
  wire 972;
  wire 973;
  wire 974;
  wire 975;
  wire 976;
  wire 977;
  wire 978;
  wire 979;
  wire 98;
  wire 980;
  wire 981;
  wire 982;
  wire 983;
  wire 984;
  wire 985;
  wire 986;
  wire 987;
  wire 988;
  wire 989;
  wire 99;
  wire 990;
  wire 991;
  wire 992;
  wire 993;
  wire 994;
  wire 995;
  wire 996;
  wire 997;
  wire 998;
  wire 999;
  wire tie_lo_T0Y0__R2_CONB_0;
  wire tie_lo_T0Y10__R2_CONB_0;
  wire tie_lo_T0Y11__R2_CONB_0;
  wire tie_lo_T0Y12__R2_CONB_0;
  wire tie_lo_T0Y13__R2_CONB_0;
  wire tie_lo_T0Y14__R2_CONB_0;
  wire tie_lo_T0Y15__R2_CONB_0;
  wire tie_lo_T0Y16__R2_CONB_0;
  wire tie_lo_T0Y17__R2_CONB_0;
  wire tie_lo_T0Y18__R2_CONB_0;
  wire tie_lo_T0Y19__R2_CONB_0;
  wire tie_lo_T0Y1__R2_CONB_0;
  wire tie_lo_T0Y20__R2_CONB_0;
  wire tie_lo_T0Y21__R2_CONB_0;
  wire tie_lo_T0Y22__R2_CONB_0;
  wire tie_lo_T0Y23__R2_CONB_0;
  wire tie_lo_T0Y24__R2_CONB_0;
  wire tie_lo_T0Y25__R2_CONB_0;
  wire tie_lo_T0Y26__R2_CONB_0;
  wire tie_lo_T0Y27__R2_CONB_0;
  wire tie_lo_T0Y28__R2_CONB_0;
  wire tie_lo_T0Y29__R2_CONB_0;
  wire tie_lo_T0Y2__R2_CONB_0;
  wire tie_lo_T0Y30__R2_CONB_0;
  wire tie_lo_T0Y31__R2_CONB_0;
  wire tie_lo_T0Y32__R2_CONB_0;
  wire tie_lo_T0Y33__R2_CONB_0;
  wire tie_lo_T0Y34__R2_CONB_0;
  wire tie_lo_T0Y35__R2_CONB_0;
  wire tie_lo_T0Y36__R2_CONB_0;
  wire tie_lo_T0Y37__R2_CONB_0;
  wire tie_lo_T0Y38__R2_CONB_0;
  wire tie_lo_T0Y39__R2_CONB_0;
  wire tie_lo_T0Y3__R2_CONB_0;
  wire tie_lo_T0Y40__R2_CONB_0;
  wire tie_lo_T0Y41__R2_CONB_0;
  wire tie_lo_T0Y42__R2_CONB_0;
  wire tie_lo_T0Y43__R2_CONB_0;
  wire tie_lo_T0Y44__R2_CONB_0;
  wire tie_lo_T0Y45__R2_CONB_0;
  wire tie_lo_T0Y46__R2_CONB_0;
  wire tie_lo_T0Y47__R2_CONB_0;
  wire tie_lo_T0Y48__R2_CONB_0;
  wire tie_lo_T0Y49__R2_CONB_0;
  wire tie_lo_T0Y4__R2_CONB_0;
  wire tie_lo_T0Y50__R2_CONB_0;
  wire tie_lo_T0Y51__R2_CONB_0;
  wire tie_lo_T0Y52__R2_CONB_0;
  wire tie_lo_T0Y53__R2_CONB_0;
  wire tie_lo_T0Y54__R2_CONB_0;
  wire tie_lo_T0Y55__R2_CONB_0;
  wire tie_lo_T0Y56__R2_CONB_0;
  wire tie_lo_T0Y57__R2_CONB_0;
  wire tie_lo_T0Y58__R2_CONB_0;
  wire tie_lo_T0Y59__R2_CONB_0;
  wire tie_lo_T0Y5__R2_CONB_0;
  wire tie_lo_T0Y60__R2_CONB_0;
  wire tie_lo_T0Y61__R2_CONB_0;
  wire tie_lo_T0Y62__R2_CONB_0;
  wire tie_lo_T0Y63__R2_CONB_0;
  wire tie_lo_T0Y64__R2_CONB_0;
  wire tie_lo_T0Y65__R2_CONB_0;
  wire tie_lo_T0Y66__R2_CONB_0;
  wire tie_lo_T0Y67__R2_CONB_0;
  wire tie_lo_T0Y68__R2_CONB_0;
  wire tie_lo_T0Y69__R2_CONB_0;
  wire tie_lo_T0Y6__R2_CONB_0;
  wire tie_lo_T0Y70__R2_CONB_0;
  wire tie_lo_T0Y71__R2_CONB_0;
  wire tie_lo_T0Y72__R2_CONB_0;
  wire tie_lo_T0Y73__R2_CONB_0;
  wire tie_lo_T0Y74__R2_CONB_0;
  wire tie_lo_T0Y75__R2_CONB_0;
  wire tie_lo_T0Y76__R2_CONB_0;
  wire tie_lo_T0Y77__R2_CONB_0;
  wire tie_lo_T0Y78__R2_CONB_0;
  wire tie_lo_T0Y79__R2_CONB_0;
  wire tie_lo_T0Y7__R2_CONB_0;
  wire tie_lo_T0Y80__R2_CONB_0;
  wire tie_lo_T0Y81__R2_CONB_0;
  wire tie_lo_T0Y82__R2_CONB_0;
  wire tie_lo_T0Y83__R2_CONB_0;
  wire tie_lo_T0Y84__R2_CONB_0;
  wire tie_lo_T0Y85__R2_CONB_0;
  wire tie_lo_T0Y86__R2_CONB_0;
  wire tie_lo_T0Y87__R2_CONB_0;
  wire tie_lo_T0Y88__R2_CONB_0;
  wire tie_lo_T0Y89__R2_CONB_0;
  wire tie_lo_T0Y8__R2_CONB_0;
  wire tie_lo_T0Y9__R2_CONB_0;
  wire tie_lo_T10Y0__R2_CONB_0;
  wire tie_lo_T10Y10__R2_CONB_0;
  wire tie_lo_T10Y11__R2_CONB_0;
  wire tie_lo_T10Y12__R2_CONB_0;
  wire tie_lo_T10Y13__R2_CONB_0;
  wire tie_lo_T10Y14__R2_CONB_0;
  wire tie_lo_T10Y15__R2_CONB_0;
  wire tie_lo_T10Y16__R2_CONB_0;
  wire tie_lo_T10Y17__R2_CONB_0;
  wire tie_lo_T10Y18__R2_CONB_0;
  wire tie_lo_T10Y19__R2_CONB_0;
  wire tie_lo_T10Y1__R2_CONB_0;
  wire tie_lo_T10Y20__R2_CONB_0;
  wire tie_lo_T10Y21__R2_CONB_0;
  wire tie_lo_T10Y22__R2_CONB_0;
  wire tie_lo_T10Y23__R2_CONB_0;
  wire tie_lo_T10Y24__R2_CONB_0;
  wire tie_lo_T10Y25__R2_CONB_0;
  wire tie_lo_T10Y26__R2_CONB_0;
  wire tie_lo_T10Y27__R2_CONB_0;
  wire tie_lo_T10Y28__R2_CONB_0;
  wire tie_lo_T10Y29__R2_CONB_0;
  wire tie_lo_T10Y2__R2_CONB_0;
  wire tie_lo_T10Y30__R2_CONB_0;
  wire tie_lo_T10Y31__R2_CONB_0;
  wire tie_lo_T10Y32__R2_CONB_0;
  wire tie_lo_T10Y33__R2_CONB_0;
  wire tie_lo_T10Y34__R2_CONB_0;
  wire tie_lo_T10Y35__R2_CONB_0;
  wire tie_lo_T10Y36__R2_CONB_0;
  wire tie_lo_T10Y37__R2_CONB_0;
  wire tie_lo_T10Y38__R2_CONB_0;
  wire tie_lo_T10Y39__R2_CONB_0;
  wire tie_lo_T10Y3__R2_CONB_0;
  wire tie_lo_T10Y40__R2_CONB_0;
  wire tie_lo_T10Y41__R2_CONB_0;
  wire tie_lo_T10Y42__R2_CONB_0;
  wire tie_lo_T10Y43__R2_CONB_0;
  wire tie_lo_T10Y44__R2_CONB_0;
  wire tie_lo_T10Y45__R2_CONB_0;
  wire tie_lo_T10Y46__R2_CONB_0;
  wire tie_lo_T10Y47__R2_CONB_0;
  wire tie_lo_T10Y48__R2_CONB_0;
  wire tie_lo_T10Y49__R2_CONB_0;
  wire tie_lo_T10Y4__R2_CONB_0;
  wire tie_lo_T10Y50__R2_CONB_0;
  wire tie_lo_T10Y51__R2_CONB_0;
  wire tie_lo_T10Y52__R2_CONB_0;
  wire tie_lo_T10Y53__R2_CONB_0;
  wire tie_lo_T10Y54__R2_CONB_0;
  wire tie_lo_T10Y55__R2_CONB_0;
  wire tie_lo_T10Y56__R2_CONB_0;
  wire tie_lo_T10Y57__R2_CONB_0;
  wire tie_lo_T10Y58__R2_CONB_0;
  wire tie_lo_T10Y59__R2_CONB_0;
  wire tie_lo_T10Y5__R2_CONB_0;
  wire tie_lo_T10Y60__R2_CONB_0;
  wire tie_lo_T10Y61__R2_CONB_0;
  wire tie_lo_T10Y62__R2_CONB_0;
  wire tie_lo_T10Y63__R2_CONB_0;
  wire tie_lo_T10Y64__R2_CONB_0;
  wire tie_lo_T10Y65__R2_CONB_0;
  wire tie_lo_T10Y66__R2_CONB_0;
  wire tie_lo_T10Y67__R2_CONB_0;
  wire tie_lo_T10Y68__R2_CONB_0;
  wire tie_lo_T10Y69__R2_CONB_0;
  wire tie_lo_T10Y6__R2_CONB_0;
  wire tie_lo_T10Y70__R2_CONB_0;
  wire tie_lo_T10Y71__R2_CONB_0;
  wire tie_lo_T10Y72__R2_CONB_0;
  wire tie_lo_T10Y73__R2_CONB_0;
  wire tie_lo_T10Y74__R2_CONB_0;
  wire tie_lo_T10Y75__R2_CONB_0;
  wire tie_lo_T10Y76__R2_CONB_0;
  wire tie_lo_T10Y77__R2_CONB_0;
  wire tie_lo_T10Y78__R2_CONB_0;
  wire tie_lo_T10Y79__R2_CONB_0;
  wire tie_lo_T10Y7__R2_CONB_0;
  wire tie_lo_T10Y80__R2_CONB_0;
  wire tie_lo_T10Y81__R2_CONB_0;
  wire tie_lo_T10Y82__R2_CONB_0;
  wire tie_lo_T10Y83__R2_CONB_0;
  wire tie_lo_T10Y84__R2_CONB_0;
  wire tie_lo_T10Y85__R2_CONB_0;
  wire tie_lo_T10Y86__R2_CONB_0;
  wire tie_lo_T10Y87__R2_CONB_0;
  wire tie_lo_T10Y88__R2_CONB_0;
  wire tie_lo_T10Y89__R2_CONB_0;
  wire tie_lo_T10Y8__R2_CONB_0;
  wire tie_lo_T10Y9__R2_CONB_0;
  wire tie_lo_T11Y0__R2_CONB_0;
  wire tie_lo_T11Y10__R2_CONB_0;
  wire tie_lo_T11Y11__R2_CONB_0;
  wire tie_lo_T11Y12__R2_CONB_0;
  wire tie_lo_T11Y13__R2_CONB_0;
  wire tie_lo_T11Y14__R2_CONB_0;
  wire tie_lo_T11Y15__R2_CONB_0;
  wire tie_lo_T11Y16__R2_CONB_0;
  wire tie_lo_T11Y17__R2_CONB_0;
  wire tie_lo_T11Y18__R2_CONB_0;
  wire tie_lo_T11Y19__R2_CONB_0;
  wire tie_lo_T11Y1__R2_CONB_0;
  wire tie_lo_T11Y20__R2_CONB_0;
  wire tie_lo_T11Y21__R2_CONB_0;
  wire tie_lo_T11Y22__R2_CONB_0;
  wire tie_lo_T11Y23__R2_CONB_0;
  wire tie_lo_T11Y24__R2_CONB_0;
  wire tie_lo_T11Y25__R2_CONB_0;
  wire tie_lo_T11Y26__R2_CONB_0;
  wire tie_lo_T11Y27__R2_CONB_0;
  wire tie_lo_T11Y28__R2_CONB_0;
  wire tie_lo_T11Y29__R2_CONB_0;
  wire tie_lo_T11Y2__R2_CONB_0;
  wire tie_lo_T11Y30__R2_CONB_0;
  wire tie_lo_T11Y31__R2_CONB_0;
  wire tie_lo_T11Y32__R2_CONB_0;
  wire tie_lo_T11Y33__R2_CONB_0;
  wire tie_lo_T11Y34__R2_CONB_0;
  wire tie_lo_T11Y35__R2_CONB_0;
  wire tie_lo_T11Y36__R2_CONB_0;
  wire tie_lo_T11Y37__R2_CONB_0;
  wire tie_lo_T11Y38__R2_CONB_0;
  wire tie_lo_T11Y39__R2_CONB_0;
  wire tie_lo_T11Y3__R2_CONB_0;
  wire tie_lo_T11Y40__R2_CONB_0;
  wire tie_lo_T11Y41__R2_CONB_0;
  wire tie_lo_T11Y42__R2_CONB_0;
  wire tie_lo_T11Y43__R2_CONB_0;
  wire tie_lo_T11Y44__R2_CONB_0;
  wire tie_lo_T11Y45__R2_CONB_0;
  wire tie_lo_T11Y46__R2_CONB_0;
  wire tie_lo_T11Y47__R2_CONB_0;
  wire tie_lo_T11Y48__R2_CONB_0;
  wire tie_lo_T11Y49__R2_CONB_0;
  wire tie_lo_T11Y4__R2_CONB_0;
  wire tie_lo_T11Y50__R2_CONB_0;
  wire tie_lo_T11Y51__R2_CONB_0;
  wire tie_lo_T11Y52__R2_CONB_0;
  wire tie_lo_T11Y53__R2_CONB_0;
  wire tie_lo_T11Y54__R2_CONB_0;
  wire tie_lo_T11Y55__R2_CONB_0;
  wire tie_lo_T11Y56__R2_CONB_0;
  wire tie_lo_T11Y57__R2_CONB_0;
  wire tie_lo_T11Y58__R2_CONB_0;
  wire tie_lo_T11Y59__R2_CONB_0;
  wire tie_lo_T11Y5__R2_CONB_0;
  wire tie_lo_T11Y60__R2_CONB_0;
  wire tie_lo_T11Y61__R2_CONB_0;
  wire tie_lo_T11Y62__R2_CONB_0;
  wire tie_lo_T11Y63__R2_CONB_0;
  wire tie_lo_T11Y64__R2_CONB_0;
  wire tie_lo_T11Y65__R2_CONB_0;
  wire tie_lo_T11Y66__R2_CONB_0;
  wire tie_lo_T11Y67__R2_CONB_0;
  wire tie_lo_T11Y68__R2_CONB_0;
  wire tie_lo_T11Y69__R2_CONB_0;
  wire tie_lo_T11Y6__R2_CONB_0;
  wire tie_lo_T11Y70__R2_CONB_0;
  wire tie_lo_T11Y71__R2_CONB_0;
  wire tie_lo_T11Y72__R2_CONB_0;
  wire tie_lo_T11Y73__R2_CONB_0;
  wire tie_lo_T11Y74__R2_CONB_0;
  wire tie_lo_T11Y75__R2_CONB_0;
  wire tie_lo_T11Y76__R2_CONB_0;
  wire tie_lo_T11Y77__R2_CONB_0;
  wire tie_lo_T11Y78__R2_CONB_0;
  wire tie_lo_T11Y79__R2_CONB_0;
  wire tie_lo_T11Y7__R2_CONB_0;
  wire tie_lo_T11Y80__R2_CONB_0;
  wire tie_lo_T11Y81__R2_CONB_0;
  wire tie_lo_T11Y82__R2_CONB_0;
  wire tie_lo_T11Y83__R2_CONB_0;
  wire tie_lo_T11Y84__R2_CONB_0;
  wire tie_lo_T11Y85__R2_CONB_0;
  wire tie_lo_T11Y86__R2_CONB_0;
  wire tie_lo_T11Y87__R2_CONB_0;
  wire tie_lo_T11Y88__R2_CONB_0;
  wire tie_lo_T11Y89__R2_CONB_0;
  wire tie_lo_T11Y8__R2_CONB_0;
  wire tie_lo_T11Y9__R2_CONB_0;
  wire tie_lo_T12Y0__R2_CONB_0;
  wire tie_lo_T12Y10__R2_CONB_0;
  wire tie_lo_T12Y11__R2_CONB_0;
  wire tie_lo_T12Y12__R2_CONB_0;
  wire tie_lo_T12Y13__R2_CONB_0;
  wire tie_lo_T12Y14__R2_CONB_0;
  wire tie_lo_T12Y15__R2_CONB_0;
  wire tie_lo_T12Y16__R2_CONB_0;
  wire tie_lo_T12Y17__R2_CONB_0;
  wire tie_lo_T12Y18__R2_CONB_0;
  wire tie_lo_T12Y19__R2_CONB_0;
  wire tie_lo_T12Y1__R2_CONB_0;
  wire tie_lo_T12Y20__R2_CONB_0;
  wire tie_lo_T12Y21__R2_CONB_0;
  wire tie_lo_T12Y22__R2_CONB_0;
  wire tie_lo_T12Y23__R2_CONB_0;
  wire tie_lo_T12Y24__R2_CONB_0;
  wire tie_lo_T12Y25__R2_CONB_0;
  wire tie_lo_T12Y26__R2_CONB_0;
  wire tie_lo_T12Y27__R2_CONB_0;
  wire tie_lo_T12Y28__R2_CONB_0;
  wire tie_lo_T12Y29__R2_CONB_0;
  wire tie_lo_T12Y2__R2_CONB_0;
  wire tie_lo_T12Y30__R2_CONB_0;
  wire tie_lo_T12Y31__R2_CONB_0;
  wire tie_lo_T12Y32__R2_CONB_0;
  wire tie_lo_T12Y33__R2_CONB_0;
  wire tie_lo_T12Y34__R2_CONB_0;
  wire tie_lo_T12Y35__R2_CONB_0;
  wire tie_lo_T12Y36__R2_CONB_0;
  wire tie_lo_T12Y37__R2_CONB_0;
  wire tie_lo_T12Y38__R2_CONB_0;
  wire tie_lo_T12Y39__R2_CONB_0;
  wire tie_lo_T12Y3__R2_CONB_0;
  wire tie_lo_T12Y40__R2_CONB_0;
  wire tie_lo_T12Y41__R2_CONB_0;
  wire tie_lo_T12Y42__R2_CONB_0;
  wire tie_lo_T12Y43__R2_CONB_0;
  wire tie_lo_T12Y44__R2_CONB_0;
  wire tie_lo_T12Y45__R2_CONB_0;
  wire tie_lo_T12Y46__R2_CONB_0;
  wire tie_lo_T12Y47__R2_CONB_0;
  wire tie_lo_T12Y48__R2_CONB_0;
  wire tie_lo_T12Y49__R2_CONB_0;
  wire tie_lo_T12Y4__R2_CONB_0;
  wire tie_lo_T12Y50__R2_CONB_0;
  wire tie_lo_T12Y51__R2_CONB_0;
  wire tie_lo_T12Y52__R2_CONB_0;
  wire tie_lo_T12Y53__R2_CONB_0;
  wire tie_lo_T12Y54__R2_CONB_0;
  wire tie_lo_T12Y55__R2_CONB_0;
  wire tie_lo_T12Y56__R2_CONB_0;
  wire tie_lo_T12Y57__R2_CONB_0;
  wire tie_lo_T12Y58__R2_CONB_0;
  wire tie_lo_T12Y59__R2_CONB_0;
  wire tie_lo_T12Y5__R2_CONB_0;
  wire tie_lo_T12Y60__R2_CONB_0;
  wire tie_lo_T12Y61__R2_CONB_0;
  wire tie_lo_T12Y62__R2_CONB_0;
  wire tie_lo_T12Y63__R2_CONB_0;
  wire tie_lo_T12Y64__R2_CONB_0;
  wire tie_lo_T12Y65__R2_CONB_0;
  wire tie_lo_T12Y66__R2_CONB_0;
  wire tie_lo_T12Y67__R2_CONB_0;
  wire tie_lo_T12Y68__R2_CONB_0;
  wire tie_lo_T12Y69__R2_CONB_0;
  wire tie_lo_T12Y6__R2_CONB_0;
  wire tie_lo_T12Y70__R2_CONB_0;
  wire tie_lo_T12Y71__R2_CONB_0;
  wire tie_lo_T12Y72__R2_CONB_0;
  wire tie_lo_T12Y73__R2_CONB_0;
  wire tie_lo_T12Y74__R2_CONB_0;
  wire tie_lo_T12Y75__R2_CONB_0;
  wire tie_lo_T12Y76__R2_CONB_0;
  wire tie_lo_T12Y77__R2_CONB_0;
  wire tie_lo_T12Y78__R2_CONB_0;
  wire tie_lo_T12Y79__R2_CONB_0;
  wire tie_lo_T12Y7__R2_CONB_0;
  wire tie_lo_T12Y80__R2_CONB_0;
  wire tie_lo_T12Y81__R2_CONB_0;
  wire tie_lo_T12Y82__R2_CONB_0;
  wire tie_lo_T12Y83__R2_CONB_0;
  wire tie_lo_T12Y84__R2_CONB_0;
  wire tie_lo_T12Y85__R2_CONB_0;
  wire tie_lo_T12Y86__R2_CONB_0;
  wire tie_lo_T12Y87__R2_CONB_0;
  wire tie_lo_T12Y88__R2_CONB_0;
  wire tie_lo_T12Y89__R2_CONB_0;
  wire tie_lo_T12Y8__R2_CONB_0;
  wire tie_lo_T12Y9__R2_CONB_0;
  wire tie_lo_T13Y0__R2_CONB_0;
  wire tie_lo_T13Y10__R2_CONB_0;
  wire tie_lo_T13Y11__R2_CONB_0;
  wire tie_lo_T13Y12__R2_CONB_0;
  wire tie_lo_T13Y13__R2_CONB_0;
  wire tie_lo_T13Y14__R2_CONB_0;
  wire tie_lo_T13Y15__R2_CONB_0;
  wire tie_lo_T13Y16__R2_CONB_0;
  wire tie_lo_T13Y17__R2_CONB_0;
  wire tie_lo_T13Y18__R2_CONB_0;
  wire tie_lo_T13Y19__R2_CONB_0;
  wire tie_lo_T13Y1__R2_CONB_0;
  wire tie_lo_T13Y20__R2_CONB_0;
  wire tie_lo_T13Y21__R2_CONB_0;
  wire tie_lo_T13Y22__R2_CONB_0;
  wire tie_lo_T13Y23__R2_CONB_0;
  wire tie_lo_T13Y24__R2_CONB_0;
  wire tie_lo_T13Y25__R2_CONB_0;
  wire tie_lo_T13Y26__R2_CONB_0;
  wire tie_lo_T13Y27__R2_CONB_0;
  wire tie_lo_T13Y28__R2_CONB_0;
  wire tie_lo_T13Y29__R2_CONB_0;
  wire tie_lo_T13Y2__R2_CONB_0;
  wire tie_lo_T13Y30__R2_CONB_0;
  wire tie_lo_T13Y31__R2_CONB_0;
  wire tie_lo_T13Y32__R2_CONB_0;
  wire tie_lo_T13Y33__R2_CONB_0;
  wire tie_lo_T13Y34__R2_CONB_0;
  wire tie_lo_T13Y35__R2_CONB_0;
  wire tie_lo_T13Y36__R2_CONB_0;
  wire tie_lo_T13Y37__R2_CONB_0;
  wire tie_lo_T13Y38__R2_CONB_0;
  wire tie_lo_T13Y39__R2_CONB_0;
  wire tie_lo_T13Y3__R2_CONB_0;
  wire tie_lo_T13Y40__R2_CONB_0;
  wire tie_lo_T13Y41__R2_CONB_0;
  wire tie_lo_T13Y42__R2_CONB_0;
  wire tie_lo_T13Y43__R2_CONB_0;
  wire tie_lo_T13Y44__R2_CONB_0;
  wire tie_lo_T13Y45__R2_CONB_0;
  wire tie_lo_T13Y46__R2_CONB_0;
  wire tie_lo_T13Y47__R2_CONB_0;
  wire tie_lo_T13Y48__R2_CONB_0;
  wire tie_lo_T13Y49__R2_CONB_0;
  wire tie_lo_T13Y4__R2_CONB_0;
  wire tie_lo_T13Y50__R2_CONB_0;
  wire tie_lo_T13Y51__R2_CONB_0;
  wire tie_lo_T13Y52__R2_CONB_0;
  wire tie_lo_T13Y53__R2_CONB_0;
  wire tie_lo_T13Y54__R2_CONB_0;
  wire tie_lo_T13Y55__R2_CONB_0;
  wire tie_lo_T13Y56__R2_CONB_0;
  wire tie_lo_T13Y57__R2_CONB_0;
  wire tie_lo_T13Y58__R2_CONB_0;
  wire tie_lo_T13Y59__R2_CONB_0;
  wire tie_lo_T13Y5__R2_CONB_0;
  wire tie_lo_T13Y60__R2_CONB_0;
  wire tie_lo_T13Y61__R2_CONB_0;
  wire tie_lo_T13Y62__R2_CONB_0;
  wire tie_lo_T13Y63__R2_CONB_0;
  wire tie_lo_T13Y64__R2_CONB_0;
  wire tie_lo_T13Y65__R2_CONB_0;
  wire tie_lo_T13Y66__R2_CONB_0;
  wire tie_lo_T13Y67__R2_CONB_0;
  wire tie_lo_T13Y68__R2_CONB_0;
  wire tie_lo_T13Y69__R2_CONB_0;
  wire tie_lo_T13Y6__R2_CONB_0;
  wire tie_lo_T13Y70__R2_CONB_0;
  wire tie_lo_T13Y71__R2_CONB_0;
  wire tie_lo_T13Y72__R2_CONB_0;
  wire tie_lo_T13Y73__R2_CONB_0;
  wire tie_lo_T13Y74__R2_CONB_0;
  wire tie_lo_T13Y75__R2_CONB_0;
  wire tie_lo_T13Y76__R2_CONB_0;
  wire tie_lo_T13Y77__R2_CONB_0;
  wire tie_lo_T13Y78__R2_CONB_0;
  wire tie_lo_T13Y79__R2_CONB_0;
  wire tie_lo_T13Y7__R2_CONB_0;
  wire tie_lo_T13Y80__R2_CONB_0;
  wire tie_lo_T13Y81__R2_CONB_0;
  wire tie_lo_T13Y82__R2_CONB_0;
  wire tie_lo_T13Y83__R2_CONB_0;
  wire tie_lo_T13Y84__R2_CONB_0;
  wire tie_lo_T13Y85__R2_CONB_0;
  wire tie_lo_T13Y86__R2_CONB_0;
  wire tie_lo_T13Y87__R2_CONB_0;
  wire tie_lo_T13Y88__R2_CONB_0;
  wire tie_lo_T13Y89__R2_CONB_0;
  wire tie_lo_T13Y8__R2_CONB_0;
  wire tie_lo_T13Y9__R2_CONB_0;
  wire tie_lo_T14Y0__R2_CONB_0;
  wire tie_lo_T14Y10__R2_CONB_0;
  wire tie_lo_T14Y11__R2_CONB_0;
  wire tie_lo_T14Y12__R2_CONB_0;
  wire tie_lo_T14Y13__R2_CONB_0;
  wire tie_lo_T14Y14__R2_CONB_0;
  wire tie_lo_T14Y15__R2_CONB_0;
  wire tie_lo_T14Y16__R2_CONB_0;
  wire tie_lo_T14Y17__R2_CONB_0;
  wire tie_lo_T14Y18__R2_CONB_0;
  wire tie_lo_T14Y19__R2_CONB_0;
  wire tie_lo_T14Y1__R2_CONB_0;
  wire tie_lo_T14Y20__R2_CONB_0;
  wire tie_lo_T14Y21__R2_CONB_0;
  wire tie_lo_T14Y22__R2_CONB_0;
  wire tie_lo_T14Y23__R2_CONB_0;
  wire tie_lo_T14Y24__R2_CONB_0;
  wire tie_lo_T14Y25__R2_CONB_0;
  wire tie_lo_T14Y26__R2_CONB_0;
  wire tie_lo_T14Y27__R2_CONB_0;
  wire tie_lo_T14Y28__R2_CONB_0;
  wire tie_lo_T14Y29__R2_CONB_0;
  wire tie_lo_T14Y2__R2_CONB_0;
  wire tie_lo_T14Y30__R2_CONB_0;
  wire tie_lo_T14Y31__R2_CONB_0;
  wire tie_lo_T14Y32__R2_CONB_0;
  wire tie_lo_T14Y33__R2_CONB_0;
  wire tie_lo_T14Y34__R2_CONB_0;
  wire tie_lo_T14Y35__R2_CONB_0;
  wire tie_lo_T14Y36__R2_CONB_0;
  wire tie_lo_T14Y37__R2_CONB_0;
  wire tie_lo_T14Y38__R2_CONB_0;
  wire tie_lo_T14Y39__R2_CONB_0;
  wire tie_lo_T14Y3__R2_CONB_0;
  wire tie_lo_T14Y40__R2_CONB_0;
  wire tie_lo_T14Y41__R2_CONB_0;
  wire tie_lo_T14Y42__R2_CONB_0;
  wire tie_lo_T14Y43__R2_CONB_0;
  wire tie_lo_T14Y44__R2_CONB_0;
  wire tie_lo_T14Y45__R2_CONB_0;
  wire tie_lo_T14Y46__R2_CONB_0;
  wire tie_lo_T14Y47__R2_CONB_0;
  wire tie_lo_T14Y48__R2_CONB_0;
  wire tie_lo_T14Y49__R2_CONB_0;
  wire tie_lo_T14Y4__R2_CONB_0;
  wire tie_lo_T14Y50__R2_CONB_0;
  wire tie_lo_T14Y51__R2_CONB_0;
  wire tie_lo_T14Y52__R2_CONB_0;
  wire tie_lo_T14Y53__R2_CONB_0;
  wire tie_lo_T14Y54__R2_CONB_0;
  wire tie_lo_T14Y55__R2_CONB_0;
  wire tie_lo_T14Y56__R2_CONB_0;
  wire tie_lo_T14Y57__R2_CONB_0;
  wire tie_lo_T14Y58__R2_CONB_0;
  wire tie_lo_T14Y59__R2_CONB_0;
  wire tie_lo_T14Y5__R2_CONB_0;
  wire tie_lo_T14Y60__R2_CONB_0;
  wire tie_lo_T14Y61__R2_CONB_0;
  wire tie_lo_T14Y62__R2_CONB_0;
  wire tie_lo_T14Y63__R2_CONB_0;
  wire tie_lo_T14Y64__R2_CONB_0;
  wire tie_lo_T14Y65__R2_CONB_0;
  wire tie_lo_T14Y66__R2_CONB_0;
  wire tie_lo_T14Y67__R2_CONB_0;
  wire tie_lo_T14Y68__R2_CONB_0;
  wire tie_lo_T14Y69__R2_CONB_0;
  wire tie_lo_T14Y6__R2_CONB_0;
  wire tie_lo_T14Y70__R2_CONB_0;
  wire tie_lo_T14Y71__R2_CONB_0;
  wire tie_lo_T14Y72__R2_CONB_0;
  wire tie_lo_T14Y73__R2_CONB_0;
  wire tie_lo_T14Y74__R2_CONB_0;
  wire tie_lo_T14Y75__R2_CONB_0;
  wire tie_lo_T14Y76__R2_CONB_0;
  wire tie_lo_T14Y77__R2_CONB_0;
  wire tie_lo_T14Y78__R2_CONB_0;
  wire tie_lo_T14Y79__R2_CONB_0;
  wire tie_lo_T14Y7__R2_CONB_0;
  wire tie_lo_T14Y80__R2_CONB_0;
  wire tie_lo_T14Y81__R2_CONB_0;
  wire tie_lo_T14Y82__R2_CONB_0;
  wire tie_lo_T14Y83__R2_CONB_0;
  wire tie_lo_T14Y84__R2_CONB_0;
  wire tie_lo_T14Y85__R2_CONB_0;
  wire tie_lo_T14Y86__R2_CONB_0;
  wire tie_lo_T14Y87__R2_CONB_0;
  wire tie_lo_T14Y88__R2_CONB_0;
  wire tie_lo_T14Y89__R2_CONB_0;
  wire tie_lo_T14Y8__R2_CONB_0;
  wire tie_lo_T14Y9__R2_CONB_0;
  wire tie_lo_T15Y0__R2_CONB_0;
  wire tie_lo_T15Y10__R2_CONB_0;
  wire tie_lo_T15Y11__R2_CONB_0;
  wire tie_lo_T15Y12__R2_CONB_0;
  wire tie_lo_T15Y13__R2_CONB_0;
  wire tie_lo_T15Y14__R2_CONB_0;
  wire tie_lo_T15Y15__R2_CONB_0;
  wire tie_lo_T15Y16__R2_CONB_0;
  wire tie_lo_T15Y17__R2_CONB_0;
  wire tie_lo_T15Y18__R2_CONB_0;
  wire tie_lo_T15Y19__R2_CONB_0;
  wire tie_lo_T15Y1__R2_CONB_0;
  wire tie_lo_T15Y20__R2_CONB_0;
  wire tie_lo_T15Y21__R2_CONB_0;
  wire tie_lo_T15Y22__R2_CONB_0;
  wire tie_lo_T15Y23__R2_CONB_0;
  wire tie_lo_T15Y24__R2_CONB_0;
  wire tie_lo_T15Y25__R2_CONB_0;
  wire tie_lo_T15Y26__R2_CONB_0;
  wire tie_lo_T15Y27__R2_CONB_0;
  wire tie_lo_T15Y28__R2_CONB_0;
  wire tie_lo_T15Y29__R2_CONB_0;
  wire tie_lo_T15Y2__R2_CONB_0;
  wire tie_lo_T15Y30__R2_CONB_0;
  wire tie_lo_T15Y31__R2_CONB_0;
  wire tie_lo_T15Y32__R2_CONB_0;
  wire tie_lo_T15Y33__R2_CONB_0;
  wire tie_lo_T15Y34__R2_CONB_0;
  wire tie_lo_T15Y35__R2_CONB_0;
  wire tie_lo_T15Y36__R2_CONB_0;
  wire tie_lo_T15Y37__R2_CONB_0;
  wire tie_lo_T15Y38__R2_CONB_0;
  wire tie_lo_T15Y39__R2_CONB_0;
  wire tie_lo_T15Y3__R2_CONB_0;
  wire tie_lo_T15Y40__R2_CONB_0;
  wire tie_lo_T15Y41__R2_CONB_0;
  wire tie_lo_T15Y42__R2_CONB_0;
  wire tie_lo_T15Y43__R2_CONB_0;
  wire tie_lo_T15Y44__R2_CONB_0;
  wire tie_lo_T15Y45__R2_CONB_0;
  wire tie_lo_T15Y46__R2_CONB_0;
  wire tie_lo_T15Y47__R2_CONB_0;
  wire tie_lo_T15Y48__R2_CONB_0;
  wire tie_lo_T15Y49__R2_CONB_0;
  wire tie_lo_T15Y4__R2_CONB_0;
  wire tie_lo_T15Y50__R2_CONB_0;
  wire tie_lo_T15Y51__R2_CONB_0;
  wire tie_lo_T15Y52__R2_CONB_0;
  wire tie_lo_T15Y53__R2_CONB_0;
  wire tie_lo_T15Y54__R2_CONB_0;
  wire tie_lo_T15Y55__R2_CONB_0;
  wire tie_lo_T15Y56__R2_CONB_0;
  wire tie_lo_T15Y57__R2_CONB_0;
  wire tie_lo_T15Y58__R2_CONB_0;
  wire tie_lo_T15Y59__R2_CONB_0;
  wire tie_lo_T15Y5__R2_CONB_0;
  wire tie_lo_T15Y60__R2_CONB_0;
  wire tie_lo_T15Y61__R2_CONB_0;
  wire tie_lo_T15Y62__R2_CONB_0;
  wire tie_lo_T15Y63__R2_CONB_0;
  wire tie_lo_T15Y64__R2_CONB_0;
  wire tie_lo_T15Y65__R2_CONB_0;
  wire tie_lo_T15Y66__R2_CONB_0;
  wire tie_lo_T15Y67__R2_CONB_0;
  wire tie_lo_T15Y68__R2_CONB_0;
  wire tie_lo_T15Y69__R2_CONB_0;
  wire tie_lo_T15Y6__R2_CONB_0;
  wire tie_lo_T15Y70__R2_CONB_0;
  wire tie_lo_T15Y71__R2_CONB_0;
  wire tie_lo_T15Y72__R2_CONB_0;
  wire tie_lo_T15Y73__R2_CONB_0;
  wire tie_lo_T15Y74__R2_CONB_0;
  wire tie_lo_T15Y75__R2_CONB_0;
  wire tie_lo_T15Y76__R2_CONB_0;
  wire tie_lo_T15Y77__R2_CONB_0;
  wire tie_lo_T15Y78__R2_CONB_0;
  wire tie_lo_T15Y79__R2_CONB_0;
  wire tie_lo_T15Y7__R2_CONB_0;
  wire tie_lo_T15Y80__R2_CONB_0;
  wire tie_lo_T15Y81__R2_CONB_0;
  wire tie_lo_T15Y82__R2_CONB_0;
  wire tie_lo_T15Y83__R2_CONB_0;
  wire tie_lo_T15Y84__R2_CONB_0;
  wire tie_lo_T15Y85__R2_CONB_0;
  wire tie_lo_T15Y86__R2_CONB_0;
  wire tie_lo_T15Y87__R2_CONB_0;
  wire tie_lo_T15Y88__R2_CONB_0;
  wire tie_lo_T15Y89__R2_CONB_0;
  wire tie_lo_T15Y8__R2_CONB_0;
  wire tie_lo_T15Y9__R2_CONB_0;
  wire tie_lo_T16Y0__R2_CONB_0;
  wire tie_lo_T16Y10__R2_CONB_0;
  wire tie_lo_T16Y11__R2_CONB_0;
  wire tie_lo_T16Y12__R2_CONB_0;
  wire tie_lo_T16Y13__R2_CONB_0;
  wire tie_lo_T16Y14__R2_CONB_0;
  wire tie_lo_T16Y15__R2_CONB_0;
  wire tie_lo_T16Y16__R2_CONB_0;
  wire tie_lo_T16Y17__R2_CONB_0;
  wire tie_lo_T16Y18__R2_CONB_0;
  wire tie_lo_T16Y19__R2_CONB_0;
  wire tie_lo_T16Y1__R2_CONB_0;
  wire tie_lo_T16Y20__R2_CONB_0;
  wire tie_lo_T16Y21__R2_CONB_0;
  wire tie_lo_T16Y22__R2_CONB_0;
  wire tie_lo_T16Y23__R2_CONB_0;
  wire tie_lo_T16Y24__R2_CONB_0;
  wire tie_lo_T16Y25__R2_CONB_0;
  wire tie_lo_T16Y26__R2_CONB_0;
  wire tie_lo_T16Y27__R2_CONB_0;
  wire tie_lo_T16Y28__R2_CONB_0;
  wire tie_lo_T16Y29__R2_CONB_0;
  wire tie_lo_T16Y2__R2_CONB_0;
  wire tie_lo_T16Y30__R2_CONB_0;
  wire tie_lo_T16Y31__R2_CONB_0;
  wire tie_lo_T16Y32__R2_CONB_0;
  wire tie_lo_T16Y33__R2_CONB_0;
  wire tie_lo_T16Y34__R2_CONB_0;
  wire tie_lo_T16Y35__R2_CONB_0;
  wire tie_lo_T16Y36__R2_CONB_0;
  wire tie_lo_T16Y37__R2_CONB_0;
  wire tie_lo_T16Y38__R2_CONB_0;
  wire tie_lo_T16Y39__R2_CONB_0;
  wire tie_lo_T16Y3__R2_CONB_0;
  wire tie_lo_T16Y40__R2_CONB_0;
  wire tie_lo_T16Y41__R2_CONB_0;
  wire tie_lo_T16Y42__R2_CONB_0;
  wire tie_lo_T16Y43__R2_CONB_0;
  wire tie_lo_T16Y44__R2_CONB_0;
  wire tie_lo_T16Y45__R2_CONB_0;
  wire tie_lo_T16Y46__R2_CONB_0;
  wire tie_lo_T16Y47__R2_CONB_0;
  wire tie_lo_T16Y48__R2_CONB_0;
  wire tie_lo_T16Y49__R2_CONB_0;
  wire tie_lo_T16Y4__R2_CONB_0;
  wire tie_lo_T16Y50__R2_CONB_0;
  wire tie_lo_T16Y51__R2_CONB_0;
  wire tie_lo_T16Y52__R2_CONB_0;
  wire tie_lo_T16Y53__R2_CONB_0;
  wire tie_lo_T16Y54__R2_CONB_0;
  wire tie_lo_T16Y55__R2_CONB_0;
  wire tie_lo_T16Y56__R2_CONB_0;
  wire tie_lo_T16Y57__R2_CONB_0;
  wire tie_lo_T16Y58__R2_CONB_0;
  wire tie_lo_T16Y59__R2_CONB_0;
  wire tie_lo_T16Y5__R2_CONB_0;
  wire tie_lo_T16Y60__R2_CONB_0;
  wire tie_lo_T16Y61__R2_CONB_0;
  wire tie_lo_T16Y62__R2_CONB_0;
  wire tie_lo_T16Y63__R2_CONB_0;
  wire tie_lo_T16Y64__R2_CONB_0;
  wire tie_lo_T16Y65__R2_CONB_0;
  wire tie_lo_T16Y66__R2_CONB_0;
  wire tie_lo_T16Y67__R2_CONB_0;
  wire tie_lo_T16Y68__R2_CONB_0;
  wire tie_lo_T16Y69__R2_CONB_0;
  wire tie_lo_T16Y6__R2_CONB_0;
  wire tie_lo_T16Y70__R2_CONB_0;
  wire tie_lo_T16Y71__R2_CONB_0;
  wire tie_lo_T16Y72__R2_CONB_0;
  wire tie_lo_T16Y73__R2_CONB_0;
  wire tie_lo_T16Y74__R2_CONB_0;
  wire tie_lo_T16Y75__R2_CONB_0;
  wire tie_lo_T16Y76__R2_CONB_0;
  wire tie_lo_T16Y77__R2_CONB_0;
  wire tie_lo_T16Y78__R2_CONB_0;
  wire tie_lo_T16Y79__R2_CONB_0;
  wire tie_lo_T16Y7__R2_CONB_0;
  wire tie_lo_T16Y80__R2_CONB_0;
  wire tie_lo_T16Y81__R2_CONB_0;
  wire tie_lo_T16Y82__R2_CONB_0;
  wire tie_lo_T16Y83__R2_CONB_0;
  wire tie_lo_T16Y84__R2_CONB_0;
  wire tie_lo_T16Y85__R2_CONB_0;
  wire tie_lo_T16Y86__R2_CONB_0;
  wire tie_lo_T16Y87__R2_CONB_0;
  wire tie_lo_T16Y88__R2_CONB_0;
  wire tie_lo_T16Y89__R2_CONB_0;
  wire tie_lo_T16Y8__R2_CONB_0;
  wire tie_lo_T16Y9__R2_CONB_0;
  wire tie_lo_T17Y0__R2_CONB_0;
  wire tie_lo_T17Y10__R2_CONB_0;
  wire tie_lo_T17Y11__R2_CONB_0;
  wire tie_lo_T17Y12__R2_CONB_0;
  wire tie_lo_T17Y13__R2_CONB_0;
  wire tie_lo_T17Y14__R2_CONB_0;
  wire tie_lo_T17Y15__R2_CONB_0;
  wire tie_lo_T17Y16__R2_CONB_0;
  wire tie_lo_T17Y17__R2_CONB_0;
  wire tie_lo_T17Y18__R2_CONB_0;
  wire tie_lo_T17Y19__R2_CONB_0;
  wire tie_lo_T17Y1__R2_CONB_0;
  wire tie_lo_T17Y20__R2_CONB_0;
  wire tie_lo_T17Y21__R2_CONB_0;
  wire tie_lo_T17Y22__R2_CONB_0;
  wire tie_lo_T17Y23__R2_CONB_0;
  wire tie_lo_T17Y24__R2_CONB_0;
  wire tie_lo_T17Y25__R2_CONB_0;
  wire tie_lo_T17Y26__R2_CONB_0;
  wire tie_lo_T17Y27__R2_CONB_0;
  wire tie_lo_T17Y28__R2_CONB_0;
  wire tie_lo_T17Y29__R2_CONB_0;
  wire tie_lo_T17Y2__R2_CONB_0;
  wire tie_lo_T17Y30__R2_CONB_0;
  wire tie_lo_T17Y31__R2_CONB_0;
  wire tie_lo_T17Y32__R2_CONB_0;
  wire tie_lo_T17Y33__R2_CONB_0;
  wire tie_lo_T17Y34__R2_CONB_0;
  wire tie_lo_T17Y35__R2_CONB_0;
  wire tie_lo_T17Y36__R2_CONB_0;
  wire tie_lo_T17Y37__R2_CONB_0;
  wire tie_lo_T17Y38__R2_CONB_0;
  wire tie_lo_T17Y39__R2_CONB_0;
  wire tie_lo_T17Y3__R2_CONB_0;
  wire tie_lo_T17Y40__R2_CONB_0;
  wire tie_lo_T17Y41__R2_CONB_0;
  wire tie_lo_T17Y42__R2_CONB_0;
  wire tie_lo_T17Y43__R2_CONB_0;
  wire tie_lo_T17Y44__R2_CONB_0;
  wire tie_lo_T17Y45__R2_CONB_0;
  wire tie_lo_T17Y46__R2_CONB_0;
  wire tie_lo_T17Y47__R2_CONB_0;
  wire tie_lo_T17Y48__R2_CONB_0;
  wire tie_lo_T17Y49__R2_CONB_0;
  wire tie_lo_T17Y4__R2_CONB_0;
  wire tie_lo_T17Y50__R2_CONB_0;
  wire tie_lo_T17Y51__R2_CONB_0;
  wire tie_lo_T17Y52__R2_CONB_0;
  wire tie_lo_T17Y53__R2_CONB_0;
  wire tie_lo_T17Y54__R2_CONB_0;
  wire tie_lo_T17Y55__R2_CONB_0;
  wire tie_lo_T17Y56__R2_CONB_0;
  wire tie_lo_T17Y57__R2_CONB_0;
  wire tie_lo_T17Y58__R2_CONB_0;
  wire tie_lo_T17Y59__R2_CONB_0;
  wire tie_lo_T17Y5__R2_CONB_0;
  wire tie_lo_T17Y60__R2_CONB_0;
  wire tie_lo_T17Y61__R2_CONB_0;
  wire tie_lo_T17Y62__R2_CONB_0;
  wire tie_lo_T17Y63__R2_CONB_0;
  wire tie_lo_T17Y64__R2_CONB_0;
  wire tie_lo_T17Y65__R2_CONB_0;
  wire tie_lo_T17Y66__R2_CONB_0;
  wire tie_lo_T17Y67__R2_CONB_0;
  wire tie_lo_T17Y68__R2_CONB_0;
  wire tie_lo_T17Y69__R2_CONB_0;
  wire tie_lo_T17Y6__R2_CONB_0;
  wire tie_lo_T17Y70__R2_CONB_0;
  wire tie_lo_T17Y71__R2_CONB_0;
  wire tie_lo_T17Y72__R2_CONB_0;
  wire tie_lo_T17Y73__R2_CONB_0;
  wire tie_lo_T17Y74__R2_CONB_0;
  wire tie_lo_T17Y75__R2_CONB_0;
  wire tie_lo_T17Y76__R2_CONB_0;
  wire tie_lo_T17Y77__R2_CONB_0;
  wire tie_lo_T17Y78__R2_CONB_0;
  wire tie_lo_T17Y79__R2_CONB_0;
  wire tie_lo_T17Y7__R2_CONB_0;
  wire tie_lo_T17Y80__R2_CONB_0;
  wire tie_lo_T17Y81__R2_CONB_0;
  wire tie_lo_T17Y82__R2_CONB_0;
  wire tie_lo_T17Y83__R2_CONB_0;
  wire tie_lo_T17Y84__R2_CONB_0;
  wire tie_lo_T17Y85__R2_CONB_0;
  wire tie_lo_T17Y86__R2_CONB_0;
  wire tie_lo_T17Y87__R2_CONB_0;
  wire tie_lo_T17Y88__R2_CONB_0;
  wire tie_lo_T17Y89__R2_CONB_0;
  wire tie_lo_T17Y8__R2_CONB_0;
  wire tie_lo_T17Y9__R2_CONB_0;
  wire tie_lo_T18Y0__R2_CONB_0;
  wire tie_lo_T18Y10__R2_CONB_0;
  wire tie_lo_T18Y11__R2_CONB_0;
  wire tie_lo_T18Y12__R2_CONB_0;
  wire tie_lo_T18Y13__R2_CONB_0;
  wire tie_lo_T18Y14__R2_CONB_0;
  wire tie_lo_T18Y15__R2_CONB_0;
  wire tie_lo_T18Y16__R2_CONB_0;
  wire tie_lo_T18Y17__R2_CONB_0;
  wire tie_lo_T18Y18__R2_CONB_0;
  wire tie_lo_T18Y19__R2_CONB_0;
  wire tie_lo_T18Y1__R2_CONB_0;
  wire tie_lo_T18Y20__R2_CONB_0;
  wire tie_lo_T18Y21__R2_CONB_0;
  wire tie_lo_T18Y22__R2_CONB_0;
  wire tie_lo_T18Y23__R2_CONB_0;
  wire tie_lo_T18Y24__R2_CONB_0;
  wire tie_lo_T18Y25__R2_CONB_0;
  wire tie_lo_T18Y26__R2_CONB_0;
  wire tie_lo_T18Y27__R2_CONB_0;
  wire tie_lo_T18Y28__R2_CONB_0;
  wire tie_lo_T18Y29__R2_CONB_0;
  wire tie_lo_T18Y2__R2_CONB_0;
  wire tie_lo_T18Y30__R2_CONB_0;
  wire tie_lo_T18Y31__R2_CONB_0;
  wire tie_lo_T18Y32__R2_CONB_0;
  wire tie_lo_T18Y33__R2_CONB_0;
  wire tie_lo_T18Y34__R2_CONB_0;
  wire tie_lo_T18Y35__R2_CONB_0;
  wire tie_lo_T18Y36__R2_CONB_0;
  wire tie_lo_T18Y37__R2_CONB_0;
  wire tie_lo_T18Y38__R2_CONB_0;
  wire tie_lo_T18Y39__R2_CONB_0;
  wire tie_lo_T18Y3__R2_CONB_0;
  wire tie_lo_T18Y40__R2_CONB_0;
  wire tie_lo_T18Y41__R2_CONB_0;
  wire tie_lo_T18Y42__R2_CONB_0;
  wire tie_lo_T18Y43__R2_CONB_0;
  wire tie_lo_T18Y44__R2_CONB_0;
  wire tie_lo_T18Y45__R2_CONB_0;
  wire tie_lo_T18Y46__R2_CONB_0;
  wire tie_lo_T18Y47__R2_CONB_0;
  wire tie_lo_T18Y48__R2_CONB_0;
  wire tie_lo_T18Y49__R2_CONB_0;
  wire tie_lo_T18Y4__R2_CONB_0;
  wire tie_lo_T18Y50__R2_CONB_0;
  wire tie_lo_T18Y51__R2_CONB_0;
  wire tie_lo_T18Y52__R2_CONB_0;
  wire tie_lo_T18Y53__R2_CONB_0;
  wire tie_lo_T18Y54__R2_CONB_0;
  wire tie_lo_T18Y55__R2_CONB_0;
  wire tie_lo_T18Y56__R2_CONB_0;
  wire tie_lo_T18Y57__R2_CONB_0;
  wire tie_lo_T18Y58__R2_CONB_0;
  wire tie_lo_T18Y59__R2_CONB_0;
  wire tie_lo_T18Y5__R2_CONB_0;
  wire tie_lo_T18Y60__R2_CONB_0;
  wire tie_lo_T18Y61__R2_CONB_0;
  wire tie_lo_T18Y62__R2_CONB_0;
  wire tie_lo_T18Y63__R2_CONB_0;
  wire tie_lo_T18Y64__R2_CONB_0;
  wire tie_lo_T18Y65__R2_CONB_0;
  wire tie_lo_T18Y66__R2_CONB_0;
  wire tie_lo_T18Y67__R2_CONB_0;
  wire tie_lo_T18Y68__R2_CONB_0;
  wire tie_lo_T18Y69__R2_CONB_0;
  wire tie_lo_T18Y6__R2_CONB_0;
  wire tie_lo_T18Y70__R2_CONB_0;
  wire tie_lo_T18Y71__R2_CONB_0;
  wire tie_lo_T18Y72__R2_CONB_0;
  wire tie_lo_T18Y73__R2_CONB_0;
  wire tie_lo_T18Y74__R2_CONB_0;
  wire tie_lo_T18Y75__R2_CONB_0;
  wire tie_lo_T18Y76__R2_CONB_0;
  wire tie_lo_T18Y77__R2_CONB_0;
  wire tie_lo_T18Y78__R2_CONB_0;
  wire tie_lo_T18Y79__R2_CONB_0;
  wire tie_lo_T18Y7__R2_CONB_0;
  wire tie_lo_T18Y80__R2_CONB_0;
  wire tie_lo_T18Y81__R2_CONB_0;
  wire tie_lo_T18Y82__R2_CONB_0;
  wire tie_lo_T18Y83__R2_CONB_0;
  wire tie_lo_T18Y84__R2_CONB_0;
  wire tie_lo_T18Y85__R2_CONB_0;
  wire tie_lo_T18Y86__R2_CONB_0;
  wire tie_lo_T18Y87__R2_CONB_0;
  wire tie_lo_T18Y88__R2_CONB_0;
  wire tie_lo_T18Y89__R2_CONB_0;
  wire tie_lo_T18Y8__R2_CONB_0;
  wire tie_lo_T18Y9__R2_CONB_0;
  wire tie_lo_T19Y0__R2_CONB_0;
  wire tie_lo_T19Y10__R2_CONB_0;
  wire tie_lo_T19Y11__R2_CONB_0;
  wire tie_lo_T19Y12__R2_CONB_0;
  wire tie_lo_T19Y13__R2_CONB_0;
  wire tie_lo_T19Y14__R2_CONB_0;
  wire tie_lo_T19Y15__R2_CONB_0;
  wire tie_lo_T19Y16__R2_CONB_0;
  wire tie_lo_T19Y17__R2_CONB_0;
  wire tie_lo_T19Y18__R2_CONB_0;
  wire tie_lo_T19Y19__R2_CONB_0;
  wire tie_lo_T19Y1__R2_CONB_0;
  wire tie_lo_T19Y20__R2_CONB_0;
  wire tie_lo_T19Y21__R2_CONB_0;
  wire tie_lo_T19Y22__R2_CONB_0;
  wire tie_lo_T19Y23__R2_CONB_0;
  wire tie_lo_T19Y24__R2_CONB_0;
  wire tie_lo_T19Y25__R2_CONB_0;
  wire tie_lo_T19Y26__R2_CONB_0;
  wire tie_lo_T19Y27__R2_CONB_0;
  wire tie_lo_T19Y28__R2_CONB_0;
  wire tie_lo_T19Y29__R2_CONB_0;
  wire tie_lo_T19Y2__R2_CONB_0;
  wire tie_lo_T19Y30__R2_CONB_0;
  wire tie_lo_T19Y31__R2_CONB_0;
  wire tie_lo_T19Y32__R2_CONB_0;
  wire tie_lo_T19Y33__R2_CONB_0;
  wire tie_lo_T19Y34__R2_CONB_0;
  wire tie_lo_T19Y35__R2_CONB_0;
  wire tie_lo_T19Y36__R2_CONB_0;
  wire tie_lo_T19Y37__R2_CONB_0;
  wire tie_lo_T19Y38__R2_CONB_0;
  wire tie_lo_T19Y39__R2_CONB_0;
  wire tie_lo_T19Y3__R2_CONB_0;
  wire tie_lo_T19Y40__R2_CONB_0;
  wire tie_lo_T19Y41__R2_CONB_0;
  wire tie_lo_T19Y42__R2_CONB_0;
  wire tie_lo_T19Y43__R2_CONB_0;
  wire tie_lo_T19Y44__R2_CONB_0;
  wire tie_lo_T19Y45__R2_CONB_0;
  wire tie_lo_T19Y46__R2_CONB_0;
  wire tie_lo_T19Y47__R2_CONB_0;
  wire tie_lo_T19Y48__R2_CONB_0;
  wire tie_lo_T19Y49__R2_CONB_0;
  wire tie_lo_T19Y4__R2_CONB_0;
  wire tie_lo_T19Y50__R2_CONB_0;
  wire tie_lo_T19Y51__R2_CONB_0;
  wire tie_lo_T19Y52__R2_CONB_0;
  wire tie_lo_T19Y53__R2_CONB_0;
  wire tie_lo_T19Y54__R2_CONB_0;
  wire tie_lo_T19Y55__R2_CONB_0;
  wire tie_lo_T19Y56__R2_CONB_0;
  wire tie_lo_T19Y57__R2_CONB_0;
  wire tie_lo_T19Y58__R2_CONB_0;
  wire tie_lo_T19Y59__R2_CONB_0;
  wire tie_lo_T19Y5__R2_CONB_0;
  wire tie_lo_T19Y60__R2_CONB_0;
  wire tie_lo_T19Y61__R2_CONB_0;
  wire tie_lo_T19Y62__R2_CONB_0;
  wire tie_lo_T19Y63__R2_CONB_0;
  wire tie_lo_T19Y64__R2_CONB_0;
  wire tie_lo_T19Y65__R2_CONB_0;
  wire tie_lo_T19Y66__R2_CONB_0;
  wire tie_lo_T19Y67__R2_CONB_0;
  wire tie_lo_T19Y68__R2_CONB_0;
  wire tie_lo_T19Y69__R2_CONB_0;
  wire tie_lo_T19Y6__R2_CONB_0;
  wire tie_lo_T19Y70__R2_CONB_0;
  wire tie_lo_T19Y71__R2_CONB_0;
  wire tie_lo_T19Y72__R2_CONB_0;
  wire tie_lo_T19Y73__R2_CONB_0;
  wire tie_lo_T19Y74__R2_CONB_0;
  wire tie_lo_T19Y75__R2_CONB_0;
  wire tie_lo_T19Y76__R2_CONB_0;
  wire tie_lo_T19Y77__R2_CONB_0;
  wire tie_lo_T19Y78__R2_CONB_0;
  wire tie_lo_T19Y79__R2_CONB_0;
  wire tie_lo_T19Y7__R2_CONB_0;
  wire tie_lo_T19Y80__R2_CONB_0;
  wire tie_lo_T19Y81__R2_CONB_0;
  wire tie_lo_T19Y82__R2_CONB_0;
  wire tie_lo_T19Y83__R2_CONB_0;
  wire tie_lo_T19Y84__R2_CONB_0;
  wire tie_lo_T19Y85__R2_CONB_0;
  wire tie_lo_T19Y86__R2_CONB_0;
  wire tie_lo_T19Y87__R2_CONB_0;
  wire tie_lo_T19Y88__R2_CONB_0;
  wire tie_lo_T19Y89__R2_CONB_0;
  wire tie_lo_T19Y8__R2_CONB_0;
  wire tie_lo_T19Y9__R2_CONB_0;
  wire tie_lo_T1Y0__R2_CONB_0;
  wire tie_lo_T1Y10__R2_CONB_0;
  wire tie_lo_T1Y11__R2_CONB_0;
  wire tie_lo_T1Y12__R2_CONB_0;
  wire tie_lo_T1Y13__R2_CONB_0;
  wire tie_lo_T1Y14__R2_CONB_0;
  wire tie_lo_T1Y15__R2_CONB_0;
  wire tie_lo_T1Y16__R2_CONB_0;
  wire tie_lo_T1Y17__R2_CONB_0;
  wire tie_lo_T1Y18__R2_CONB_0;
  wire tie_lo_T1Y19__R2_CONB_0;
  wire tie_lo_T1Y1__R2_CONB_0;
  wire tie_lo_T1Y20__R2_CONB_0;
  wire tie_lo_T1Y21__R2_CONB_0;
  wire tie_lo_T1Y22__R2_CONB_0;
  wire tie_lo_T1Y23__R2_CONB_0;
  wire tie_lo_T1Y24__R2_CONB_0;
  wire tie_lo_T1Y25__R2_CONB_0;
  wire tie_lo_T1Y26__R2_CONB_0;
  wire tie_lo_T1Y27__R2_CONB_0;
  wire tie_lo_T1Y28__R2_CONB_0;
  wire tie_lo_T1Y29__R2_CONB_0;
  wire tie_lo_T1Y2__R2_CONB_0;
  wire tie_lo_T1Y30__R2_CONB_0;
  wire tie_lo_T1Y31__R2_CONB_0;
  wire tie_lo_T1Y32__R2_CONB_0;
  wire tie_lo_T1Y33__R2_CONB_0;
  wire tie_lo_T1Y34__R2_CONB_0;
  wire tie_lo_T1Y35__R2_CONB_0;
  wire tie_lo_T1Y36__R2_CONB_0;
  wire tie_lo_T1Y37__R2_CONB_0;
  wire tie_lo_T1Y38__R2_CONB_0;
  wire tie_lo_T1Y39__R2_CONB_0;
  wire tie_lo_T1Y3__R2_CONB_0;
  wire tie_lo_T1Y40__R2_CONB_0;
  wire tie_lo_T1Y41__R2_CONB_0;
  wire tie_lo_T1Y42__R2_CONB_0;
  wire tie_lo_T1Y43__R2_CONB_0;
  wire tie_lo_T1Y44__R2_CONB_0;
  wire tie_lo_T1Y45__R2_CONB_0;
  wire tie_lo_T1Y46__R2_CONB_0;
  wire tie_lo_T1Y47__R2_CONB_0;
  wire tie_lo_T1Y48__R2_CONB_0;
  wire tie_lo_T1Y49__R2_CONB_0;
  wire tie_lo_T1Y4__R2_CONB_0;
  wire tie_lo_T1Y50__R2_CONB_0;
  wire tie_lo_T1Y51__R2_CONB_0;
  wire tie_lo_T1Y52__R2_CONB_0;
  wire tie_lo_T1Y53__R2_CONB_0;
  wire tie_lo_T1Y54__R2_CONB_0;
  wire tie_lo_T1Y55__R2_CONB_0;
  wire tie_lo_T1Y56__R2_CONB_0;
  wire tie_lo_T1Y57__R2_CONB_0;
  wire tie_lo_T1Y58__R2_CONB_0;
  wire tie_lo_T1Y59__R2_CONB_0;
  wire tie_lo_T1Y5__R2_CONB_0;
  wire tie_lo_T1Y60__R2_CONB_0;
  wire tie_lo_T1Y61__R2_CONB_0;
  wire tie_lo_T1Y62__R2_CONB_0;
  wire tie_lo_T1Y63__R2_CONB_0;
  wire tie_lo_T1Y64__R2_CONB_0;
  wire tie_lo_T1Y65__R2_CONB_0;
  wire tie_lo_T1Y66__R2_CONB_0;
  wire tie_lo_T1Y67__R2_CONB_0;
  wire tie_lo_T1Y68__R2_CONB_0;
  wire tie_lo_T1Y69__R2_CONB_0;
  wire tie_lo_T1Y6__R2_CONB_0;
  wire tie_lo_T1Y70__R2_CONB_0;
  wire tie_lo_T1Y71__R2_CONB_0;
  wire tie_lo_T1Y72__R2_CONB_0;
  wire tie_lo_T1Y73__R2_CONB_0;
  wire tie_lo_T1Y74__R2_CONB_0;
  wire tie_lo_T1Y75__R2_CONB_0;
  wire tie_lo_T1Y76__R2_CONB_0;
  wire tie_lo_T1Y77__R2_CONB_0;
  wire tie_lo_T1Y78__R2_CONB_0;
  wire tie_lo_T1Y79__R2_CONB_0;
  wire tie_lo_T1Y7__R2_CONB_0;
  wire tie_lo_T1Y80__R2_CONB_0;
  wire tie_lo_T1Y81__R2_CONB_0;
  wire tie_lo_T1Y82__R2_CONB_0;
  wire tie_lo_T1Y83__R2_CONB_0;
  wire tie_lo_T1Y84__R2_CONB_0;
  wire tie_lo_T1Y85__R2_CONB_0;
  wire tie_lo_T1Y86__R2_CONB_0;
  wire tie_lo_T1Y87__R2_CONB_0;
  wire tie_lo_T1Y88__R2_CONB_0;
  wire tie_lo_T1Y89__R2_CONB_0;
  wire tie_lo_T1Y8__R2_CONB_0;
  wire tie_lo_T1Y9__R2_CONB_0;
  wire tie_lo_T20Y0__R2_CONB_0;
  wire tie_lo_T20Y10__R2_CONB_0;
  wire tie_lo_T20Y11__R2_CONB_0;
  wire tie_lo_T20Y12__R2_CONB_0;
  wire tie_lo_T20Y13__R2_CONB_0;
  wire tie_lo_T20Y14__R2_CONB_0;
  wire tie_lo_T20Y15__R2_CONB_0;
  wire tie_lo_T20Y16__R2_CONB_0;
  wire tie_lo_T20Y17__R2_CONB_0;
  wire tie_lo_T20Y18__R2_CONB_0;
  wire tie_lo_T20Y19__R2_CONB_0;
  wire tie_lo_T20Y1__R2_CONB_0;
  wire tie_lo_T20Y20__R2_CONB_0;
  wire tie_lo_T20Y21__R2_CONB_0;
  wire tie_lo_T20Y22__R2_CONB_0;
  wire tie_lo_T20Y23__R2_CONB_0;
  wire tie_lo_T20Y24__R2_CONB_0;
  wire tie_lo_T20Y25__R2_CONB_0;
  wire tie_lo_T20Y26__R2_CONB_0;
  wire tie_lo_T20Y27__R2_CONB_0;
  wire tie_lo_T20Y28__R2_CONB_0;
  wire tie_lo_T20Y29__R2_CONB_0;
  wire tie_lo_T20Y2__R2_CONB_0;
  wire tie_lo_T20Y30__R2_CONB_0;
  wire tie_lo_T20Y31__R2_CONB_0;
  wire tie_lo_T20Y32__R2_CONB_0;
  wire tie_lo_T20Y33__R2_CONB_0;
  wire tie_lo_T20Y34__R2_CONB_0;
  wire tie_lo_T20Y35__R2_CONB_0;
  wire tie_lo_T20Y36__R2_CONB_0;
  wire tie_lo_T20Y37__R2_CONB_0;
  wire tie_lo_T20Y38__R2_CONB_0;
  wire tie_lo_T20Y39__R2_CONB_0;
  wire tie_lo_T20Y3__R2_CONB_0;
  wire tie_lo_T20Y40__R2_CONB_0;
  wire tie_lo_T20Y41__R2_CONB_0;
  wire tie_lo_T20Y42__R2_CONB_0;
  wire tie_lo_T20Y43__R2_CONB_0;
  wire tie_lo_T20Y44__R2_CONB_0;
  wire tie_lo_T20Y45__R2_CONB_0;
  wire tie_lo_T20Y46__R2_CONB_0;
  wire tie_lo_T20Y47__R2_CONB_0;
  wire tie_lo_T20Y48__R2_CONB_0;
  wire tie_lo_T20Y49__R2_CONB_0;
  wire tie_lo_T20Y4__R2_CONB_0;
  wire tie_lo_T20Y50__R2_CONB_0;
  wire tie_lo_T20Y51__R2_CONB_0;
  wire tie_lo_T20Y52__R2_CONB_0;
  wire tie_lo_T20Y53__R2_CONB_0;
  wire tie_lo_T20Y54__R2_CONB_0;
  wire tie_lo_T20Y55__R2_CONB_0;
  wire tie_lo_T20Y56__R2_CONB_0;
  wire tie_lo_T20Y57__R2_CONB_0;
  wire tie_lo_T20Y58__R2_CONB_0;
  wire tie_lo_T20Y59__R2_CONB_0;
  wire tie_lo_T20Y5__R2_CONB_0;
  wire tie_lo_T20Y60__R2_CONB_0;
  wire tie_lo_T20Y61__R2_CONB_0;
  wire tie_lo_T20Y62__R2_CONB_0;
  wire tie_lo_T20Y63__R2_CONB_0;
  wire tie_lo_T20Y64__R2_CONB_0;
  wire tie_lo_T20Y65__R2_CONB_0;
  wire tie_lo_T20Y66__R2_CONB_0;
  wire tie_lo_T20Y67__R2_CONB_0;
  wire tie_lo_T20Y68__R2_CONB_0;
  wire tie_lo_T20Y69__R2_CONB_0;
  wire tie_lo_T20Y6__R2_CONB_0;
  wire tie_lo_T20Y70__R2_CONB_0;
  wire tie_lo_T20Y71__R2_CONB_0;
  wire tie_lo_T20Y72__R2_CONB_0;
  wire tie_lo_T20Y73__R2_CONB_0;
  wire tie_lo_T20Y74__R2_CONB_0;
  wire tie_lo_T20Y75__R2_CONB_0;
  wire tie_lo_T20Y76__R2_CONB_0;
  wire tie_lo_T20Y77__R2_CONB_0;
  wire tie_lo_T20Y78__R2_CONB_0;
  wire tie_lo_T20Y79__R2_CONB_0;
  wire tie_lo_T20Y7__R2_CONB_0;
  wire tie_lo_T20Y80__R2_CONB_0;
  wire tie_lo_T20Y81__R2_CONB_0;
  wire tie_lo_T20Y82__R2_CONB_0;
  wire tie_lo_T20Y83__R2_CONB_0;
  wire tie_lo_T20Y84__R2_CONB_0;
  wire tie_lo_T20Y85__R2_CONB_0;
  wire tie_lo_T20Y86__R2_CONB_0;
  wire tie_lo_T20Y87__R2_CONB_0;
  wire tie_lo_T20Y88__R2_CONB_0;
  wire tie_lo_T20Y89__R2_CONB_0;
  wire tie_lo_T20Y8__R2_CONB_0;
  wire tie_lo_T20Y9__R2_CONB_0;
  wire tie_lo_T21Y0__R2_CONB_0;
  wire tie_lo_T21Y10__R2_CONB_0;
  wire tie_lo_T21Y11__R2_CONB_0;
  wire tie_lo_T21Y12__R2_CONB_0;
  wire tie_lo_T21Y13__R2_CONB_0;
  wire tie_lo_T21Y14__R2_CONB_0;
  wire tie_lo_T21Y15__R2_CONB_0;
  wire tie_lo_T21Y16__R2_CONB_0;
  wire tie_lo_T21Y17__R2_CONB_0;
  wire tie_lo_T21Y18__R2_CONB_0;
  wire tie_lo_T21Y19__R2_CONB_0;
  wire tie_lo_T21Y1__R2_CONB_0;
  wire tie_lo_T21Y20__R2_CONB_0;
  wire tie_lo_T21Y21__R2_CONB_0;
  wire tie_lo_T21Y22__R2_CONB_0;
  wire tie_lo_T21Y23__R2_CONB_0;
  wire tie_lo_T21Y24__R2_CONB_0;
  wire tie_lo_T21Y25__R2_CONB_0;
  wire tie_lo_T21Y26__R2_CONB_0;
  wire tie_lo_T21Y27__R2_CONB_0;
  wire tie_lo_T21Y28__R2_CONB_0;
  wire tie_lo_T21Y29__R2_CONB_0;
  wire tie_lo_T21Y2__R2_CONB_0;
  wire tie_lo_T21Y30__R2_CONB_0;
  wire tie_lo_T21Y31__R2_CONB_0;
  wire tie_lo_T21Y32__R2_CONB_0;
  wire tie_lo_T21Y33__R2_CONB_0;
  wire tie_lo_T21Y34__R2_CONB_0;
  wire tie_lo_T21Y35__R2_CONB_0;
  wire tie_lo_T21Y36__R2_CONB_0;
  wire tie_lo_T21Y37__R2_CONB_0;
  wire tie_lo_T21Y38__R2_CONB_0;
  wire tie_lo_T21Y39__R2_CONB_0;
  wire tie_lo_T21Y3__R2_CONB_0;
  wire tie_lo_T21Y40__R2_CONB_0;
  wire tie_lo_T21Y41__R2_CONB_0;
  wire tie_lo_T21Y42__R2_CONB_0;
  wire tie_lo_T21Y43__R2_CONB_0;
  wire tie_lo_T21Y44__R2_CONB_0;
  wire tie_lo_T21Y45__R2_CONB_0;
  wire tie_lo_T21Y46__R2_CONB_0;
  wire tie_lo_T21Y47__R2_CONB_0;
  wire tie_lo_T21Y48__R2_CONB_0;
  wire tie_lo_T21Y49__R2_CONB_0;
  wire tie_lo_T21Y4__R2_CONB_0;
  wire tie_lo_T21Y50__R2_CONB_0;
  wire tie_lo_T21Y51__R2_CONB_0;
  wire tie_lo_T21Y52__R2_CONB_0;
  wire tie_lo_T21Y53__R2_CONB_0;
  wire tie_lo_T21Y54__R2_CONB_0;
  wire tie_lo_T21Y55__R2_CONB_0;
  wire tie_lo_T21Y56__R2_CONB_0;
  wire tie_lo_T21Y57__R2_CONB_0;
  wire tie_lo_T21Y58__R2_CONB_0;
  wire tie_lo_T21Y59__R2_CONB_0;
  wire tie_lo_T21Y5__R2_CONB_0;
  wire tie_lo_T21Y60__R2_CONB_0;
  wire tie_lo_T21Y61__R2_CONB_0;
  wire tie_lo_T21Y62__R2_CONB_0;
  wire tie_lo_T21Y63__R2_CONB_0;
  wire tie_lo_T21Y64__R2_CONB_0;
  wire tie_lo_T21Y65__R2_CONB_0;
  wire tie_lo_T21Y66__R2_CONB_0;
  wire tie_lo_T21Y67__R2_CONB_0;
  wire tie_lo_T21Y68__R2_CONB_0;
  wire tie_lo_T21Y69__R2_CONB_0;
  wire tie_lo_T21Y6__R2_CONB_0;
  wire tie_lo_T21Y70__R2_CONB_0;
  wire tie_lo_T21Y71__R2_CONB_0;
  wire tie_lo_T21Y72__R2_CONB_0;
  wire tie_lo_T21Y73__R2_CONB_0;
  wire tie_lo_T21Y74__R2_CONB_0;
  wire tie_lo_T21Y75__R2_CONB_0;
  wire tie_lo_T21Y76__R2_CONB_0;
  wire tie_lo_T21Y77__R2_CONB_0;
  wire tie_lo_T21Y78__R2_CONB_0;
  wire tie_lo_T21Y79__R2_CONB_0;
  wire tie_lo_T21Y7__R2_CONB_0;
  wire tie_lo_T21Y80__R2_CONB_0;
  wire tie_lo_T21Y81__R2_CONB_0;
  wire tie_lo_T21Y82__R2_CONB_0;
  wire tie_lo_T21Y83__R2_CONB_0;
  wire tie_lo_T21Y84__R2_CONB_0;
  wire tie_lo_T21Y85__R2_CONB_0;
  wire tie_lo_T21Y86__R2_CONB_0;
  wire tie_lo_T21Y87__R2_CONB_0;
  wire tie_lo_T21Y88__R2_CONB_0;
  wire tie_lo_T21Y89__R2_CONB_0;
  wire tie_lo_T21Y8__R2_CONB_0;
  wire tie_lo_T21Y9__R2_CONB_0;
  wire tie_lo_T22Y0__R2_CONB_0;
  wire tie_lo_T22Y10__R2_CONB_0;
  wire tie_lo_T22Y11__R2_CONB_0;
  wire tie_lo_T22Y12__R2_CONB_0;
  wire tie_lo_T22Y13__R2_CONB_0;
  wire tie_lo_T22Y14__R2_CONB_0;
  wire tie_lo_T22Y15__R2_CONB_0;
  wire tie_lo_T22Y16__R2_CONB_0;
  wire tie_lo_T22Y17__R2_CONB_0;
  wire tie_lo_T22Y18__R2_CONB_0;
  wire tie_lo_T22Y19__R2_CONB_0;
  wire tie_lo_T22Y1__R2_CONB_0;
  wire tie_lo_T22Y20__R2_CONB_0;
  wire tie_lo_T22Y21__R2_CONB_0;
  wire tie_lo_T22Y22__R2_CONB_0;
  wire tie_lo_T22Y23__R2_CONB_0;
  wire tie_lo_T22Y24__R2_CONB_0;
  wire tie_lo_T22Y25__R2_CONB_0;
  wire tie_lo_T22Y26__R2_CONB_0;
  wire tie_lo_T22Y27__R2_CONB_0;
  wire tie_lo_T22Y28__R2_CONB_0;
  wire tie_lo_T22Y29__R2_CONB_0;
  wire tie_lo_T22Y2__R2_CONB_0;
  wire tie_lo_T22Y30__R2_CONB_0;
  wire tie_lo_T22Y31__R2_CONB_0;
  wire tie_lo_T22Y32__R2_CONB_0;
  wire tie_lo_T22Y33__R2_CONB_0;
  wire tie_lo_T22Y34__R2_CONB_0;
  wire tie_lo_T22Y35__R2_CONB_0;
  wire tie_lo_T22Y36__R2_CONB_0;
  wire tie_lo_T22Y37__R2_CONB_0;
  wire tie_lo_T22Y38__R2_CONB_0;
  wire tie_lo_T22Y39__R2_CONB_0;
  wire tie_lo_T22Y3__R2_CONB_0;
  wire tie_lo_T22Y40__R2_CONB_0;
  wire tie_lo_T22Y41__R2_CONB_0;
  wire tie_lo_T22Y42__R2_CONB_0;
  wire tie_lo_T22Y43__R2_CONB_0;
  wire tie_lo_T22Y44__R2_CONB_0;
  wire tie_lo_T22Y45__R2_CONB_0;
  wire tie_lo_T22Y46__R2_CONB_0;
  wire tie_lo_T22Y47__R2_CONB_0;
  wire tie_lo_T22Y48__R2_CONB_0;
  wire tie_lo_T22Y49__R2_CONB_0;
  wire tie_lo_T22Y4__R2_CONB_0;
  wire tie_lo_T22Y50__R2_CONB_0;
  wire tie_lo_T22Y51__R2_CONB_0;
  wire tie_lo_T22Y52__R2_CONB_0;
  wire tie_lo_T22Y53__R2_CONB_0;
  wire tie_lo_T22Y54__R2_CONB_0;
  wire tie_lo_T22Y55__R2_CONB_0;
  wire tie_lo_T22Y56__R2_CONB_0;
  wire tie_lo_T22Y57__R2_CONB_0;
  wire tie_lo_T22Y58__R2_CONB_0;
  wire tie_lo_T22Y59__R2_CONB_0;
  wire tie_lo_T22Y5__R2_CONB_0;
  wire tie_lo_T22Y60__R2_CONB_0;
  wire tie_lo_T22Y61__R2_CONB_0;
  wire tie_lo_T22Y62__R2_CONB_0;
  wire tie_lo_T22Y63__R2_CONB_0;
  wire tie_lo_T22Y64__R2_CONB_0;
  wire tie_lo_T22Y65__R2_CONB_0;
  wire tie_lo_T22Y66__R2_CONB_0;
  wire tie_lo_T22Y67__R2_CONB_0;
  wire tie_lo_T22Y68__R2_CONB_0;
  wire tie_lo_T22Y69__R2_CONB_0;
  wire tie_lo_T22Y6__R2_CONB_0;
  wire tie_lo_T22Y70__R2_CONB_0;
  wire tie_lo_T22Y71__R2_CONB_0;
  wire tie_lo_T22Y72__R2_CONB_0;
  wire tie_lo_T22Y73__R2_CONB_0;
  wire tie_lo_T22Y74__R2_CONB_0;
  wire tie_lo_T22Y75__R2_CONB_0;
  wire tie_lo_T22Y76__R2_CONB_0;
  wire tie_lo_T22Y77__R2_CONB_0;
  wire tie_lo_T22Y78__R2_CONB_0;
  wire tie_lo_T22Y79__R2_CONB_0;
  wire tie_lo_T22Y7__R2_CONB_0;
  wire tie_lo_T22Y80__R2_CONB_0;
  wire tie_lo_T22Y81__R2_CONB_0;
  wire tie_lo_T22Y82__R2_CONB_0;
  wire tie_lo_T22Y83__R2_CONB_0;
  wire tie_lo_T22Y84__R2_CONB_0;
  wire tie_lo_T22Y85__R2_CONB_0;
  wire tie_lo_T22Y86__R2_CONB_0;
  wire tie_lo_T22Y87__R2_CONB_0;
  wire tie_lo_T22Y88__R2_CONB_0;
  wire tie_lo_T22Y89__R2_CONB_0;
  wire tie_lo_T22Y8__R2_CONB_0;
  wire tie_lo_T22Y9__R2_CONB_0;
  wire tie_lo_T23Y0__R2_CONB_0;
  wire tie_lo_T23Y10__R2_CONB_0;
  wire tie_lo_T23Y11__R2_CONB_0;
  wire tie_lo_T23Y12__R2_CONB_0;
  wire tie_lo_T23Y13__R2_CONB_0;
  wire tie_lo_T23Y14__R2_CONB_0;
  wire tie_lo_T23Y15__R2_CONB_0;
  wire tie_lo_T23Y16__R2_CONB_0;
  wire tie_lo_T23Y17__R2_CONB_0;
  wire tie_lo_T23Y18__R2_CONB_0;
  wire tie_lo_T23Y19__R2_CONB_0;
  wire tie_lo_T23Y1__R2_CONB_0;
  wire tie_lo_T23Y20__R2_CONB_0;
  wire tie_lo_T23Y21__R2_CONB_0;
  wire tie_lo_T23Y22__R2_CONB_0;
  wire tie_lo_T23Y23__R2_CONB_0;
  wire tie_lo_T23Y24__R2_CONB_0;
  wire tie_lo_T23Y25__R2_CONB_0;
  wire tie_lo_T23Y26__R2_CONB_0;
  wire tie_lo_T23Y27__R2_CONB_0;
  wire tie_lo_T23Y28__R2_CONB_0;
  wire tie_lo_T23Y29__R2_CONB_0;
  wire tie_lo_T23Y2__R2_CONB_0;
  wire tie_lo_T23Y30__R2_CONB_0;
  wire tie_lo_T23Y31__R2_CONB_0;
  wire tie_lo_T23Y32__R2_CONB_0;
  wire tie_lo_T23Y33__R2_CONB_0;
  wire tie_lo_T23Y34__R2_CONB_0;
  wire tie_lo_T23Y35__R2_CONB_0;
  wire tie_lo_T23Y36__R2_CONB_0;
  wire tie_lo_T23Y37__R2_CONB_0;
  wire tie_lo_T23Y38__R2_CONB_0;
  wire tie_lo_T23Y39__R2_CONB_0;
  wire tie_lo_T23Y3__R2_CONB_0;
  wire tie_lo_T23Y40__R2_CONB_0;
  wire tie_lo_T23Y41__R2_CONB_0;
  wire tie_lo_T23Y42__R2_CONB_0;
  wire tie_lo_T23Y43__R2_CONB_0;
  wire tie_lo_T23Y44__R2_CONB_0;
  wire tie_lo_T23Y45__R2_CONB_0;
  wire tie_lo_T23Y46__R2_CONB_0;
  wire tie_lo_T23Y47__R2_CONB_0;
  wire tie_lo_T23Y48__R2_CONB_0;
  wire tie_lo_T23Y49__R2_CONB_0;
  wire tie_lo_T23Y4__R2_CONB_0;
  wire tie_lo_T23Y50__R2_CONB_0;
  wire tie_lo_T23Y51__R2_CONB_0;
  wire tie_lo_T23Y52__R2_CONB_0;
  wire tie_lo_T23Y53__R2_CONB_0;
  wire tie_lo_T23Y54__R2_CONB_0;
  wire tie_lo_T23Y55__R2_CONB_0;
  wire tie_lo_T23Y56__R2_CONB_0;
  wire tie_lo_T23Y57__R2_CONB_0;
  wire tie_lo_T23Y58__R2_CONB_0;
  wire tie_lo_T23Y59__R2_CONB_0;
  wire tie_lo_T23Y5__R2_CONB_0;
  wire tie_lo_T23Y60__R2_CONB_0;
  wire tie_lo_T23Y61__R2_CONB_0;
  wire tie_lo_T23Y62__R2_CONB_0;
  wire tie_lo_T23Y63__R2_CONB_0;
  wire tie_lo_T23Y64__R2_CONB_0;
  wire tie_lo_T23Y65__R2_CONB_0;
  wire tie_lo_T23Y66__R2_CONB_0;
  wire tie_lo_T23Y67__R2_CONB_0;
  wire tie_lo_T23Y68__R2_CONB_0;
  wire tie_lo_T23Y69__R2_CONB_0;
  wire tie_lo_T23Y6__R2_CONB_0;
  wire tie_lo_T23Y70__R2_CONB_0;
  wire tie_lo_T23Y71__R2_CONB_0;
  wire tie_lo_T23Y72__R2_CONB_0;
  wire tie_lo_T23Y73__R2_CONB_0;
  wire tie_lo_T23Y74__R2_CONB_0;
  wire tie_lo_T23Y75__R2_CONB_0;
  wire tie_lo_T23Y76__R2_CONB_0;
  wire tie_lo_T23Y77__R2_CONB_0;
  wire tie_lo_T23Y78__R2_CONB_0;
  wire tie_lo_T23Y79__R2_CONB_0;
  wire tie_lo_T23Y7__R2_CONB_0;
  wire tie_lo_T23Y80__R2_CONB_0;
  wire tie_lo_T23Y81__R2_CONB_0;
  wire tie_lo_T23Y82__R2_CONB_0;
  wire tie_lo_T23Y83__R2_CONB_0;
  wire tie_lo_T23Y84__R2_CONB_0;
  wire tie_lo_T23Y85__R2_CONB_0;
  wire tie_lo_T23Y86__R2_CONB_0;
  wire tie_lo_T23Y87__R2_CONB_0;
  wire tie_lo_T23Y88__R2_CONB_0;
  wire tie_lo_T23Y89__R2_CONB_0;
  wire tie_lo_T23Y8__R2_CONB_0;
  wire tie_lo_T23Y9__R2_CONB_0;
  wire tie_lo_T24Y0__R2_CONB_0;
  wire tie_lo_T24Y10__R2_CONB_0;
  wire tie_lo_T24Y11__R2_CONB_0;
  wire tie_lo_T24Y12__R2_CONB_0;
  wire tie_lo_T24Y13__R2_CONB_0;
  wire tie_lo_T24Y14__R2_CONB_0;
  wire tie_lo_T24Y15__R2_CONB_0;
  wire tie_lo_T24Y16__R2_CONB_0;
  wire tie_lo_T24Y17__R2_CONB_0;
  wire tie_lo_T24Y18__R2_CONB_0;
  wire tie_lo_T24Y19__R2_CONB_0;
  wire tie_lo_T24Y1__R2_CONB_0;
  wire tie_lo_T24Y20__R2_CONB_0;
  wire tie_lo_T24Y21__R2_CONB_0;
  wire tie_lo_T24Y22__R2_CONB_0;
  wire tie_lo_T24Y23__R2_CONB_0;
  wire tie_lo_T24Y24__R2_CONB_0;
  wire tie_lo_T24Y25__R2_CONB_0;
  wire tie_lo_T24Y26__R2_CONB_0;
  wire tie_lo_T24Y27__R2_CONB_0;
  wire tie_lo_T24Y28__R2_CONB_0;
  wire tie_lo_T24Y29__R2_CONB_0;
  wire tie_lo_T24Y2__R2_CONB_0;
  wire tie_lo_T24Y30__R2_CONB_0;
  wire tie_lo_T24Y31__R2_CONB_0;
  wire tie_lo_T24Y32__R2_CONB_0;
  wire tie_lo_T24Y33__R2_CONB_0;
  wire tie_lo_T24Y34__R2_CONB_0;
  wire tie_lo_T24Y35__R2_CONB_0;
  wire tie_lo_T24Y36__R2_CONB_0;
  wire tie_lo_T24Y37__R2_CONB_0;
  wire tie_lo_T24Y38__R2_CONB_0;
  wire tie_lo_T24Y39__R2_CONB_0;
  wire tie_lo_T24Y3__R2_CONB_0;
  wire tie_lo_T24Y40__R2_CONB_0;
  wire tie_lo_T24Y41__R2_CONB_0;
  wire tie_lo_T24Y42__R2_CONB_0;
  wire tie_lo_T24Y43__R2_CONB_0;
  wire tie_lo_T24Y44__R2_CONB_0;
  wire tie_lo_T24Y45__R2_CONB_0;
  wire tie_lo_T24Y46__R2_CONB_0;
  wire tie_lo_T24Y47__R2_CONB_0;
  wire tie_lo_T24Y48__R2_CONB_0;
  wire tie_lo_T24Y49__R2_CONB_0;
  wire tie_lo_T24Y4__R2_CONB_0;
  wire tie_lo_T24Y50__R2_CONB_0;
  wire tie_lo_T24Y51__R2_CONB_0;
  wire tie_lo_T24Y52__R2_CONB_0;
  wire tie_lo_T24Y53__R2_CONB_0;
  wire tie_lo_T24Y54__R2_CONB_0;
  wire tie_lo_T24Y55__R2_CONB_0;
  wire tie_lo_T24Y56__R2_CONB_0;
  wire tie_lo_T24Y57__R2_CONB_0;
  wire tie_lo_T24Y58__R2_CONB_0;
  wire tie_lo_T24Y59__R2_CONB_0;
  wire tie_lo_T24Y5__R2_CONB_0;
  wire tie_lo_T24Y60__R2_CONB_0;
  wire tie_lo_T24Y61__R2_CONB_0;
  wire tie_lo_T24Y62__R2_CONB_0;
  wire tie_lo_T24Y63__R2_CONB_0;
  wire tie_lo_T24Y64__R2_CONB_0;
  wire tie_lo_T24Y65__R2_CONB_0;
  wire tie_lo_T24Y66__R2_CONB_0;
  wire tie_lo_T24Y67__R2_CONB_0;
  wire tie_lo_T24Y68__R2_CONB_0;
  wire tie_lo_T24Y69__R2_CONB_0;
  wire tie_lo_T24Y6__R2_CONB_0;
  wire tie_lo_T24Y70__R2_CONB_0;
  wire tie_lo_T24Y71__R2_CONB_0;
  wire tie_lo_T24Y72__R2_CONB_0;
  wire tie_lo_T24Y73__R2_CONB_0;
  wire tie_lo_T24Y74__R2_CONB_0;
  wire tie_lo_T24Y75__R2_CONB_0;
  wire tie_lo_T24Y76__R2_CONB_0;
  wire tie_lo_T24Y77__R2_CONB_0;
  wire tie_lo_T24Y78__R2_CONB_0;
  wire tie_lo_T24Y79__R2_CONB_0;
  wire tie_lo_T24Y7__R2_CONB_0;
  wire tie_lo_T24Y80__R2_CONB_0;
  wire tie_lo_T24Y81__R2_CONB_0;
  wire tie_lo_T24Y82__R2_CONB_0;
  wire tie_lo_T24Y83__R2_CONB_0;
  wire tie_lo_T24Y84__R2_CONB_0;
  wire tie_lo_T24Y85__R2_CONB_0;
  wire tie_lo_T24Y86__R2_CONB_0;
  wire tie_lo_T24Y87__R2_CONB_0;
  wire tie_lo_T24Y88__R2_CONB_0;
  wire tie_lo_T24Y89__R2_CONB_0;
  wire tie_lo_T24Y8__R2_CONB_0;
  wire tie_lo_T24Y9__R2_CONB_0;
  wire tie_lo_T25Y0__R2_CONB_0;
  wire tie_lo_T25Y10__R2_CONB_0;
  wire tie_lo_T25Y11__R2_CONB_0;
  wire tie_lo_T25Y12__R2_CONB_0;
  wire tie_lo_T25Y13__R2_CONB_0;
  wire tie_lo_T25Y14__R2_CONB_0;
  wire tie_lo_T25Y15__R2_CONB_0;
  wire tie_lo_T25Y16__R2_CONB_0;
  wire tie_lo_T25Y17__R2_CONB_0;
  wire tie_lo_T25Y18__R2_CONB_0;
  wire tie_lo_T25Y19__R2_CONB_0;
  wire tie_lo_T25Y1__R2_CONB_0;
  wire tie_lo_T25Y20__R2_CONB_0;
  wire tie_lo_T25Y21__R2_CONB_0;
  wire tie_lo_T25Y22__R2_CONB_0;
  wire tie_lo_T25Y23__R2_CONB_0;
  wire tie_lo_T25Y24__R2_CONB_0;
  wire tie_lo_T25Y25__R2_CONB_0;
  wire tie_lo_T25Y26__R2_CONB_0;
  wire tie_lo_T25Y27__R2_CONB_0;
  wire tie_lo_T25Y28__R2_CONB_0;
  wire tie_lo_T25Y29__R2_CONB_0;
  wire tie_lo_T25Y2__R2_CONB_0;
  wire tie_lo_T25Y30__R2_CONB_0;
  wire tie_lo_T25Y31__R2_CONB_0;
  wire tie_lo_T25Y32__R2_CONB_0;
  wire tie_lo_T25Y33__R2_CONB_0;
  wire tie_lo_T25Y34__R2_CONB_0;
  wire tie_lo_T25Y35__R2_CONB_0;
  wire tie_lo_T25Y36__R2_CONB_0;
  wire tie_lo_T25Y37__R2_CONB_0;
  wire tie_lo_T25Y38__R2_CONB_0;
  wire tie_lo_T25Y39__R2_CONB_0;
  wire tie_lo_T25Y3__R2_CONB_0;
  wire tie_lo_T25Y40__R2_CONB_0;
  wire tie_lo_T25Y41__R2_CONB_0;
  wire tie_lo_T25Y42__R2_CONB_0;
  wire tie_lo_T25Y43__R2_CONB_0;
  wire tie_lo_T25Y44__R2_CONB_0;
  wire tie_lo_T25Y45__R2_CONB_0;
  wire tie_lo_T25Y46__R2_CONB_0;
  wire tie_lo_T25Y47__R2_CONB_0;
  wire tie_lo_T25Y48__R2_CONB_0;
  wire tie_lo_T25Y49__R2_CONB_0;
  wire tie_lo_T25Y4__R2_CONB_0;
  wire tie_lo_T25Y50__R2_CONB_0;
  wire tie_lo_T25Y51__R2_CONB_0;
  wire tie_lo_T25Y52__R2_CONB_0;
  wire tie_lo_T25Y53__R2_CONB_0;
  wire tie_lo_T25Y54__R2_CONB_0;
  wire tie_lo_T25Y55__R2_CONB_0;
  wire tie_lo_T25Y56__R2_CONB_0;
  wire tie_lo_T25Y57__R2_CONB_0;
  wire tie_lo_T25Y58__R2_CONB_0;
  wire tie_lo_T25Y59__R2_CONB_0;
  wire tie_lo_T25Y5__R2_CONB_0;
  wire tie_lo_T25Y60__R2_CONB_0;
  wire tie_lo_T25Y61__R2_CONB_0;
  wire tie_lo_T25Y62__R2_CONB_0;
  wire tie_lo_T25Y63__R2_CONB_0;
  wire tie_lo_T25Y64__R2_CONB_0;
  wire tie_lo_T25Y65__R2_CONB_0;
  wire tie_lo_T25Y66__R2_CONB_0;
  wire tie_lo_T25Y67__R2_CONB_0;
  wire tie_lo_T25Y68__R2_CONB_0;
  wire tie_lo_T25Y69__R2_CONB_0;
  wire tie_lo_T25Y6__R2_CONB_0;
  wire tie_lo_T25Y70__R2_CONB_0;
  wire tie_lo_T25Y71__R2_CONB_0;
  wire tie_lo_T25Y72__R2_CONB_0;
  wire tie_lo_T25Y73__R2_CONB_0;
  wire tie_lo_T25Y74__R2_CONB_0;
  wire tie_lo_T25Y75__R2_CONB_0;
  wire tie_lo_T25Y76__R2_CONB_0;
  wire tie_lo_T25Y77__R2_CONB_0;
  wire tie_lo_T25Y78__R2_CONB_0;
  wire tie_lo_T25Y79__R2_CONB_0;
  wire tie_lo_T25Y7__R2_CONB_0;
  wire tie_lo_T25Y80__R2_CONB_0;
  wire tie_lo_T25Y81__R2_CONB_0;
  wire tie_lo_T25Y82__R2_CONB_0;
  wire tie_lo_T25Y83__R2_CONB_0;
  wire tie_lo_T25Y84__R2_CONB_0;
  wire tie_lo_T25Y85__R2_CONB_0;
  wire tie_lo_T25Y86__R2_CONB_0;
  wire tie_lo_T25Y87__R2_CONB_0;
  wire tie_lo_T25Y88__R2_CONB_0;
  wire tie_lo_T25Y89__R2_CONB_0;
  wire tie_lo_T25Y8__R2_CONB_0;
  wire tie_lo_T25Y9__R2_CONB_0;
  wire tie_lo_T26Y0__R2_CONB_0;
  wire tie_lo_T26Y10__R2_CONB_0;
  wire tie_lo_T26Y11__R2_CONB_0;
  wire tie_lo_T26Y12__R2_CONB_0;
  wire tie_lo_T26Y13__R2_CONB_0;
  wire tie_lo_T26Y14__R2_CONB_0;
  wire tie_lo_T26Y15__R2_CONB_0;
  wire tie_lo_T26Y16__R2_CONB_0;
  wire tie_lo_T26Y17__R2_CONB_0;
  wire tie_lo_T26Y18__R2_CONB_0;
  wire tie_lo_T26Y19__R2_CONB_0;
  wire tie_lo_T26Y1__R2_CONB_0;
  wire tie_lo_T26Y20__R2_CONB_0;
  wire tie_lo_T26Y21__R2_CONB_0;
  wire tie_lo_T26Y22__R2_CONB_0;
  wire tie_lo_T26Y23__R2_CONB_0;
  wire tie_lo_T26Y24__R2_CONB_0;
  wire tie_lo_T26Y25__R2_CONB_0;
  wire tie_lo_T26Y26__R2_CONB_0;
  wire tie_lo_T26Y27__R2_CONB_0;
  wire tie_lo_T26Y28__R2_CONB_0;
  wire tie_lo_T26Y29__R2_CONB_0;
  wire tie_lo_T26Y2__R2_CONB_0;
  wire tie_lo_T26Y30__R2_CONB_0;
  wire tie_lo_T26Y31__R2_CONB_0;
  wire tie_lo_T26Y32__R2_CONB_0;
  wire tie_lo_T26Y33__R2_CONB_0;
  wire tie_lo_T26Y34__R2_CONB_0;
  wire tie_lo_T26Y35__R2_CONB_0;
  wire tie_lo_T26Y36__R2_CONB_0;
  wire tie_lo_T26Y37__R2_CONB_0;
  wire tie_lo_T26Y38__R2_CONB_0;
  wire tie_lo_T26Y39__R2_CONB_0;
  wire tie_lo_T26Y3__R2_CONB_0;
  wire tie_lo_T26Y40__R2_CONB_0;
  wire tie_lo_T26Y41__R2_CONB_0;
  wire tie_lo_T26Y42__R2_CONB_0;
  wire tie_lo_T26Y43__R2_CONB_0;
  wire tie_lo_T26Y44__R2_CONB_0;
  wire tie_lo_T26Y45__R2_CONB_0;
  wire tie_lo_T26Y46__R2_CONB_0;
  wire tie_lo_T26Y47__R2_CONB_0;
  wire tie_lo_T26Y48__R2_CONB_0;
  wire tie_lo_T26Y49__R2_CONB_0;
  wire tie_lo_T26Y4__R2_CONB_0;
  wire tie_lo_T26Y50__R2_CONB_0;
  wire tie_lo_T26Y51__R2_CONB_0;
  wire tie_lo_T26Y52__R2_CONB_0;
  wire tie_lo_T26Y53__R2_CONB_0;
  wire tie_lo_T26Y54__R2_CONB_0;
  wire tie_lo_T26Y55__R2_CONB_0;
  wire tie_lo_T26Y56__R2_CONB_0;
  wire tie_lo_T26Y57__R2_CONB_0;
  wire tie_lo_T26Y58__R2_CONB_0;
  wire tie_lo_T26Y59__R2_CONB_0;
  wire tie_lo_T26Y5__R2_CONB_0;
  wire tie_lo_T26Y60__R2_CONB_0;
  wire tie_lo_T26Y61__R2_CONB_0;
  wire tie_lo_T26Y62__R2_CONB_0;
  wire tie_lo_T26Y63__R2_CONB_0;
  wire tie_lo_T26Y64__R2_CONB_0;
  wire tie_lo_T26Y65__R2_CONB_0;
  wire tie_lo_T26Y66__R2_CONB_0;
  wire tie_lo_T26Y67__R2_CONB_0;
  wire tie_lo_T26Y68__R2_CONB_0;
  wire tie_lo_T26Y69__R2_CONB_0;
  wire tie_lo_T26Y6__R2_CONB_0;
  wire tie_lo_T26Y70__R2_CONB_0;
  wire tie_lo_T26Y71__R2_CONB_0;
  wire tie_lo_T26Y72__R2_CONB_0;
  wire tie_lo_T26Y73__R2_CONB_0;
  wire tie_lo_T26Y74__R2_CONB_0;
  wire tie_lo_T26Y75__R2_CONB_0;
  wire tie_lo_T26Y76__R2_CONB_0;
  wire tie_lo_T26Y77__R2_CONB_0;
  wire tie_lo_T26Y78__R2_CONB_0;
  wire tie_lo_T26Y79__R2_CONB_0;
  wire tie_lo_T26Y7__R2_CONB_0;
  wire tie_lo_T26Y80__R2_CONB_0;
  wire tie_lo_T26Y81__R2_CONB_0;
  wire tie_lo_T26Y82__R2_CONB_0;
  wire tie_lo_T26Y83__R2_CONB_0;
  wire tie_lo_T26Y84__R2_CONB_0;
  wire tie_lo_T26Y85__R2_CONB_0;
  wire tie_lo_T26Y86__R2_CONB_0;
  wire tie_lo_T26Y87__R2_CONB_0;
  wire tie_lo_T26Y88__R2_CONB_0;
  wire tie_lo_T26Y89__R2_CONB_0;
  wire tie_lo_T26Y8__R2_CONB_0;
  wire tie_lo_T26Y9__R2_CONB_0;
  wire tie_lo_T27Y0__R2_CONB_0;
  wire tie_lo_T27Y10__R2_CONB_0;
  wire tie_lo_T27Y11__R2_CONB_0;
  wire tie_lo_T27Y12__R2_CONB_0;
  wire tie_lo_T27Y13__R2_CONB_0;
  wire tie_lo_T27Y14__R2_CONB_0;
  wire tie_lo_T27Y15__R2_CONB_0;
  wire tie_lo_T27Y16__R2_CONB_0;
  wire tie_lo_T27Y17__R2_CONB_0;
  wire tie_lo_T27Y18__R2_CONB_0;
  wire tie_lo_T27Y19__R2_CONB_0;
  wire tie_lo_T27Y1__R2_CONB_0;
  wire tie_lo_T27Y20__R2_CONB_0;
  wire tie_lo_T27Y21__R2_CONB_0;
  wire tie_lo_T27Y22__R2_CONB_0;
  wire tie_lo_T27Y23__R2_CONB_0;
  wire tie_lo_T27Y24__R2_CONB_0;
  wire tie_lo_T27Y25__R2_CONB_0;
  wire tie_lo_T27Y26__R2_CONB_0;
  wire tie_lo_T27Y27__R2_CONB_0;
  wire tie_lo_T27Y28__R2_CONB_0;
  wire tie_lo_T27Y29__R2_CONB_0;
  wire tie_lo_T27Y2__R2_CONB_0;
  wire tie_lo_T27Y30__R2_CONB_0;
  wire tie_lo_T27Y31__R2_CONB_0;
  wire tie_lo_T27Y32__R2_CONB_0;
  wire tie_lo_T27Y33__R2_CONB_0;
  wire tie_lo_T27Y34__R2_CONB_0;
  wire tie_lo_T27Y35__R2_CONB_0;
  wire tie_lo_T27Y36__R2_CONB_0;
  wire tie_lo_T27Y37__R2_CONB_0;
  wire tie_lo_T27Y38__R2_CONB_0;
  wire tie_lo_T27Y39__R2_CONB_0;
  wire tie_lo_T27Y3__R2_CONB_0;
  wire tie_lo_T27Y40__R2_CONB_0;
  wire tie_lo_T27Y41__R2_CONB_0;
  wire tie_lo_T27Y42__R2_CONB_0;
  wire tie_lo_T27Y43__R2_CONB_0;
  wire tie_lo_T27Y44__R2_CONB_0;
  wire tie_lo_T27Y45__R2_CONB_0;
  wire tie_lo_T27Y46__R2_CONB_0;
  wire tie_lo_T27Y47__R2_CONB_0;
  wire tie_lo_T27Y48__R2_CONB_0;
  wire tie_lo_T27Y49__R2_CONB_0;
  wire tie_lo_T27Y4__R2_CONB_0;
  wire tie_lo_T27Y50__R2_CONB_0;
  wire tie_lo_T27Y51__R2_CONB_0;
  wire tie_lo_T27Y52__R2_CONB_0;
  wire tie_lo_T27Y53__R2_CONB_0;
  wire tie_lo_T27Y54__R2_CONB_0;
  wire tie_lo_T27Y55__R2_CONB_0;
  wire tie_lo_T27Y56__R2_CONB_0;
  wire tie_lo_T27Y57__R2_CONB_0;
  wire tie_lo_T27Y58__R2_CONB_0;
  wire tie_lo_T27Y59__R2_CONB_0;
  wire tie_lo_T27Y5__R2_CONB_0;
  wire tie_lo_T27Y60__R2_CONB_0;
  wire tie_lo_T27Y61__R2_CONB_0;
  wire tie_lo_T27Y62__R2_CONB_0;
  wire tie_lo_T27Y63__R2_CONB_0;
  wire tie_lo_T27Y64__R2_CONB_0;
  wire tie_lo_T27Y65__R2_CONB_0;
  wire tie_lo_T27Y66__R2_CONB_0;
  wire tie_lo_T27Y67__R2_CONB_0;
  wire tie_lo_T27Y68__R2_CONB_0;
  wire tie_lo_T27Y69__R2_CONB_0;
  wire tie_lo_T27Y6__R2_CONB_0;
  wire tie_lo_T27Y70__R2_CONB_0;
  wire tie_lo_T27Y71__R2_CONB_0;
  wire tie_lo_T27Y72__R2_CONB_0;
  wire tie_lo_T27Y73__R2_CONB_0;
  wire tie_lo_T27Y74__R2_CONB_0;
  wire tie_lo_T27Y75__R2_CONB_0;
  wire tie_lo_T27Y76__R2_CONB_0;
  wire tie_lo_T27Y77__R2_CONB_0;
  wire tie_lo_T27Y78__R2_CONB_0;
  wire tie_lo_T27Y79__R2_CONB_0;
  wire tie_lo_T27Y7__R2_CONB_0;
  wire tie_lo_T27Y80__R2_CONB_0;
  wire tie_lo_T27Y81__R2_CONB_0;
  wire tie_lo_T27Y82__R2_CONB_0;
  wire tie_lo_T27Y83__R2_CONB_0;
  wire tie_lo_T27Y84__R2_CONB_0;
  wire tie_lo_T27Y85__R2_CONB_0;
  wire tie_lo_T27Y86__R2_CONB_0;
  wire tie_lo_T27Y87__R2_CONB_0;
  wire tie_lo_T27Y88__R2_CONB_0;
  wire tie_lo_T27Y89__R2_CONB_0;
  wire tie_lo_T27Y8__R2_CONB_0;
  wire tie_lo_T27Y9__R2_CONB_0;
  wire tie_lo_T28Y0__R2_CONB_0;
  wire tie_lo_T28Y10__R2_CONB_0;
  wire tie_lo_T28Y11__R2_CONB_0;
  wire tie_lo_T28Y12__R2_CONB_0;
  wire tie_lo_T28Y13__R2_CONB_0;
  wire tie_lo_T28Y14__R2_CONB_0;
  wire tie_lo_T28Y15__R2_CONB_0;
  wire tie_lo_T28Y16__R2_CONB_0;
  wire tie_lo_T28Y17__R2_CONB_0;
  wire tie_lo_T28Y18__R2_CONB_0;
  wire tie_lo_T28Y19__R2_CONB_0;
  wire tie_lo_T28Y1__R2_CONB_0;
  wire tie_lo_T28Y20__R2_CONB_0;
  wire tie_lo_T28Y21__R2_CONB_0;
  wire tie_lo_T28Y22__R2_CONB_0;
  wire tie_lo_T28Y23__R2_CONB_0;
  wire tie_lo_T28Y24__R2_CONB_0;
  wire tie_lo_T28Y25__R2_CONB_0;
  wire tie_lo_T28Y26__R2_CONB_0;
  wire tie_lo_T28Y27__R2_CONB_0;
  wire tie_lo_T28Y28__R2_CONB_0;
  wire tie_lo_T28Y29__R2_CONB_0;
  wire tie_lo_T28Y2__R2_CONB_0;
  wire tie_lo_T28Y30__R2_CONB_0;
  wire tie_lo_T28Y31__R2_CONB_0;
  wire tie_lo_T28Y32__R2_CONB_0;
  wire tie_lo_T28Y33__R2_CONB_0;
  wire tie_lo_T28Y34__R2_CONB_0;
  wire tie_lo_T28Y35__R2_CONB_0;
  wire tie_lo_T28Y36__R2_CONB_0;
  wire tie_lo_T28Y37__R2_CONB_0;
  wire tie_lo_T28Y38__R2_CONB_0;
  wire tie_lo_T28Y39__R2_CONB_0;
  wire tie_lo_T28Y3__R2_CONB_0;
  wire tie_lo_T28Y40__R2_CONB_0;
  wire tie_lo_T28Y41__R2_CONB_0;
  wire tie_lo_T28Y42__R2_CONB_0;
  wire tie_lo_T28Y43__R2_CONB_0;
  wire tie_lo_T28Y44__R2_CONB_0;
  wire tie_lo_T28Y45__R2_CONB_0;
  wire tie_lo_T28Y46__R2_CONB_0;
  wire tie_lo_T28Y47__R2_CONB_0;
  wire tie_lo_T28Y48__R2_CONB_0;
  wire tie_lo_T28Y49__R2_CONB_0;
  wire tie_lo_T28Y4__R2_CONB_0;
  wire tie_lo_T28Y50__R2_CONB_0;
  wire tie_lo_T28Y51__R2_CONB_0;
  wire tie_lo_T28Y52__R2_CONB_0;
  wire tie_lo_T28Y53__R2_CONB_0;
  wire tie_lo_T28Y54__R2_CONB_0;
  wire tie_lo_T28Y55__R2_CONB_0;
  wire tie_lo_T28Y56__R2_CONB_0;
  wire tie_lo_T28Y57__R2_CONB_0;
  wire tie_lo_T28Y58__R2_CONB_0;
  wire tie_lo_T28Y59__R2_CONB_0;
  wire tie_lo_T28Y5__R2_CONB_0;
  wire tie_lo_T28Y60__R2_CONB_0;
  wire tie_lo_T28Y61__R2_CONB_0;
  wire tie_lo_T28Y62__R2_CONB_0;
  wire tie_lo_T28Y63__R2_CONB_0;
  wire tie_lo_T28Y64__R2_CONB_0;
  wire tie_lo_T28Y65__R2_CONB_0;
  wire tie_lo_T28Y66__R2_CONB_0;
  wire tie_lo_T28Y67__R2_CONB_0;
  wire tie_lo_T28Y68__R2_CONB_0;
  wire tie_lo_T28Y69__R2_CONB_0;
  wire tie_lo_T28Y6__R2_CONB_0;
  wire tie_lo_T28Y70__R2_CONB_0;
  wire tie_lo_T28Y71__R2_CONB_0;
  wire tie_lo_T28Y72__R2_CONB_0;
  wire tie_lo_T28Y73__R2_CONB_0;
  wire tie_lo_T28Y74__R2_CONB_0;
  wire tie_lo_T28Y75__R2_CONB_0;
  wire tie_lo_T28Y76__R2_CONB_0;
  wire tie_lo_T28Y77__R2_CONB_0;
  wire tie_lo_T28Y78__R2_CONB_0;
  wire tie_lo_T28Y79__R2_CONB_0;
  wire tie_lo_T28Y7__R2_CONB_0;
  wire tie_lo_T28Y80__R2_CONB_0;
  wire tie_lo_T28Y81__R2_CONB_0;
  wire tie_lo_T28Y82__R2_CONB_0;
  wire tie_lo_T28Y83__R2_CONB_0;
  wire tie_lo_T28Y84__R2_CONB_0;
  wire tie_lo_T28Y85__R2_CONB_0;
  wire tie_lo_T28Y86__R2_CONB_0;
  wire tie_lo_T28Y87__R2_CONB_0;
  wire tie_lo_T28Y88__R2_CONB_0;
  wire tie_lo_T28Y89__R2_CONB_0;
  wire tie_lo_T28Y8__R2_CONB_0;
  wire tie_lo_T28Y9__R2_CONB_0;
  wire tie_lo_T29Y0__R2_CONB_0;
  wire tie_lo_T29Y10__R2_CONB_0;
  wire tie_lo_T29Y11__R2_CONB_0;
  wire tie_lo_T29Y12__R2_CONB_0;
  wire tie_lo_T29Y13__R2_CONB_0;
  wire tie_lo_T29Y14__R2_CONB_0;
  wire tie_lo_T29Y15__R2_CONB_0;
  wire tie_lo_T29Y16__R2_CONB_0;
  wire tie_lo_T29Y17__R2_CONB_0;
  wire tie_lo_T29Y18__R2_CONB_0;
  wire tie_lo_T29Y19__R2_CONB_0;
  wire tie_lo_T29Y1__R2_CONB_0;
  wire tie_lo_T29Y20__R2_CONB_0;
  wire tie_lo_T29Y21__R2_CONB_0;
  wire tie_lo_T29Y22__R2_CONB_0;
  wire tie_lo_T29Y23__R2_CONB_0;
  wire tie_lo_T29Y24__R2_CONB_0;
  wire tie_lo_T29Y25__R2_CONB_0;
  wire tie_lo_T29Y26__R2_CONB_0;
  wire tie_lo_T29Y27__R2_CONB_0;
  wire tie_lo_T29Y28__R2_CONB_0;
  wire tie_lo_T29Y29__R2_CONB_0;
  wire tie_lo_T29Y2__R2_CONB_0;
  wire tie_lo_T29Y30__R2_CONB_0;
  wire tie_lo_T29Y31__R2_CONB_0;
  wire tie_lo_T29Y32__R2_CONB_0;
  wire tie_lo_T29Y33__R2_CONB_0;
  wire tie_lo_T29Y34__R2_CONB_0;
  wire tie_lo_T29Y35__R2_CONB_0;
  wire tie_lo_T29Y36__R2_CONB_0;
  wire tie_lo_T29Y37__R2_CONB_0;
  wire tie_lo_T29Y38__R2_CONB_0;
  wire tie_lo_T29Y39__R2_CONB_0;
  wire tie_lo_T29Y3__R2_CONB_0;
  wire tie_lo_T29Y40__R2_CONB_0;
  wire tie_lo_T29Y41__R2_CONB_0;
  wire tie_lo_T29Y42__R2_CONB_0;
  wire tie_lo_T29Y43__R2_CONB_0;
  wire tie_lo_T29Y44__R2_CONB_0;
  wire tie_lo_T29Y45__R2_CONB_0;
  wire tie_lo_T29Y46__R2_CONB_0;
  wire tie_lo_T29Y47__R2_CONB_0;
  wire tie_lo_T29Y48__R2_CONB_0;
  wire tie_lo_T29Y49__R2_CONB_0;
  wire tie_lo_T29Y4__R2_CONB_0;
  wire tie_lo_T29Y50__R2_CONB_0;
  wire tie_lo_T29Y51__R2_CONB_0;
  wire tie_lo_T29Y52__R2_CONB_0;
  wire tie_lo_T29Y53__R2_CONB_0;
  wire tie_lo_T29Y54__R2_CONB_0;
  wire tie_lo_T29Y55__R2_CONB_0;
  wire tie_lo_T29Y56__R2_CONB_0;
  wire tie_lo_T29Y57__R2_CONB_0;
  wire tie_lo_T29Y58__R2_CONB_0;
  wire tie_lo_T29Y59__R2_CONB_0;
  wire tie_lo_T29Y5__R2_CONB_0;
  wire tie_lo_T29Y60__R2_CONB_0;
  wire tie_lo_T29Y61__R2_CONB_0;
  wire tie_lo_T29Y62__R2_CONB_0;
  wire tie_lo_T29Y63__R2_CONB_0;
  wire tie_lo_T29Y64__R2_CONB_0;
  wire tie_lo_T29Y65__R2_CONB_0;
  wire tie_lo_T29Y66__R2_CONB_0;
  wire tie_lo_T29Y67__R2_CONB_0;
  wire tie_lo_T29Y68__R2_CONB_0;
  wire tie_lo_T29Y69__R2_CONB_0;
  wire tie_lo_T29Y6__R2_CONB_0;
  wire tie_lo_T29Y70__R2_CONB_0;
  wire tie_lo_T29Y71__R2_CONB_0;
  wire tie_lo_T29Y72__R2_CONB_0;
  wire tie_lo_T29Y73__R2_CONB_0;
  wire tie_lo_T29Y74__R2_CONB_0;
  wire tie_lo_T29Y75__R2_CONB_0;
  wire tie_lo_T29Y76__R2_CONB_0;
  wire tie_lo_T29Y77__R2_CONB_0;
  wire tie_lo_T29Y78__R2_CONB_0;
  wire tie_lo_T29Y79__R2_CONB_0;
  wire tie_lo_T29Y7__R2_CONB_0;
  wire tie_lo_T29Y80__R2_CONB_0;
  wire tie_lo_T29Y81__R2_CONB_0;
  wire tie_lo_T29Y82__R2_CONB_0;
  wire tie_lo_T29Y83__R2_CONB_0;
  wire tie_lo_T29Y84__R2_CONB_0;
  wire tie_lo_T29Y85__R2_CONB_0;
  wire tie_lo_T29Y86__R2_CONB_0;
  wire tie_lo_T29Y87__R2_CONB_0;
  wire tie_lo_T29Y88__R2_CONB_0;
  wire tie_lo_T29Y89__R2_CONB_0;
  wire tie_lo_T29Y8__R2_CONB_0;
  wire tie_lo_T29Y9__R2_CONB_0;
  wire tie_lo_T2Y0__R2_CONB_0;
  wire tie_lo_T2Y10__R2_CONB_0;
  wire tie_lo_T2Y11__R2_CONB_0;
  wire tie_lo_T2Y12__R2_CONB_0;
  wire tie_lo_T2Y13__R2_CONB_0;
  wire tie_lo_T2Y14__R2_CONB_0;
  wire tie_lo_T2Y15__R2_CONB_0;
  wire tie_lo_T2Y16__R2_CONB_0;
  wire tie_lo_T2Y17__R2_CONB_0;
  wire tie_lo_T2Y18__R2_CONB_0;
  wire tie_lo_T2Y19__R2_CONB_0;
  wire tie_lo_T2Y1__R2_CONB_0;
  wire tie_lo_T2Y20__R2_CONB_0;
  wire tie_lo_T2Y21__R2_CONB_0;
  wire tie_lo_T2Y22__R2_CONB_0;
  wire tie_lo_T2Y23__R2_CONB_0;
  wire tie_lo_T2Y24__R2_CONB_0;
  wire tie_lo_T2Y25__R2_CONB_0;
  wire tie_lo_T2Y26__R2_CONB_0;
  wire tie_lo_T2Y27__R2_CONB_0;
  wire tie_lo_T2Y28__R2_CONB_0;
  wire tie_lo_T2Y29__R2_CONB_0;
  wire tie_lo_T2Y2__R2_CONB_0;
  wire tie_lo_T2Y30__R2_CONB_0;
  wire tie_lo_T2Y31__R2_CONB_0;
  wire tie_lo_T2Y32__R2_CONB_0;
  wire tie_lo_T2Y33__R2_CONB_0;
  wire tie_lo_T2Y34__R2_CONB_0;
  wire tie_lo_T2Y35__R2_CONB_0;
  wire tie_lo_T2Y36__R2_CONB_0;
  wire tie_lo_T2Y37__R2_CONB_0;
  wire tie_lo_T2Y38__R2_CONB_0;
  wire tie_lo_T2Y39__R2_CONB_0;
  wire tie_lo_T2Y3__R2_CONB_0;
  wire tie_lo_T2Y40__R2_CONB_0;
  wire tie_lo_T2Y41__R2_CONB_0;
  wire tie_lo_T2Y42__R2_CONB_0;
  wire tie_lo_T2Y43__R2_CONB_0;
  wire tie_lo_T2Y44__R2_CONB_0;
  wire tie_lo_T2Y45__R2_CONB_0;
  wire tie_lo_T2Y46__R2_CONB_0;
  wire tie_lo_T2Y47__R2_CONB_0;
  wire tie_lo_T2Y48__R2_CONB_0;
  wire tie_lo_T2Y49__R2_CONB_0;
  wire tie_lo_T2Y4__R2_CONB_0;
  wire tie_lo_T2Y50__R2_CONB_0;
  wire tie_lo_T2Y51__R2_CONB_0;
  wire tie_lo_T2Y52__R2_CONB_0;
  wire tie_lo_T2Y53__R2_CONB_0;
  wire tie_lo_T2Y54__R2_CONB_0;
  wire tie_lo_T2Y55__R2_CONB_0;
  wire tie_lo_T2Y56__R2_CONB_0;
  wire tie_lo_T2Y57__R2_CONB_0;
  wire tie_lo_T2Y58__R2_CONB_0;
  wire tie_lo_T2Y59__R2_CONB_0;
  wire tie_lo_T2Y5__R2_CONB_0;
  wire tie_lo_T2Y60__R2_CONB_0;
  wire tie_lo_T2Y61__R2_CONB_0;
  wire tie_lo_T2Y62__R2_CONB_0;
  wire tie_lo_T2Y63__R2_CONB_0;
  wire tie_lo_T2Y64__R2_CONB_0;
  wire tie_lo_T2Y65__R2_CONB_0;
  wire tie_lo_T2Y66__R2_CONB_0;
  wire tie_lo_T2Y67__R2_CONB_0;
  wire tie_lo_T2Y68__R2_CONB_0;
  wire tie_lo_T2Y69__R2_CONB_0;
  wire tie_lo_T2Y6__R2_CONB_0;
  wire tie_lo_T2Y70__R2_CONB_0;
  wire tie_lo_T2Y71__R2_CONB_0;
  wire tie_lo_T2Y72__R2_CONB_0;
  wire tie_lo_T2Y73__R2_CONB_0;
  wire tie_lo_T2Y74__R2_CONB_0;
  wire tie_lo_T2Y75__R2_CONB_0;
  wire tie_lo_T2Y76__R2_CONB_0;
  wire tie_lo_T2Y77__R2_CONB_0;
  wire tie_lo_T2Y78__R2_CONB_0;
  wire tie_lo_T2Y79__R2_CONB_0;
  wire tie_lo_T2Y7__R2_CONB_0;
  wire tie_lo_T2Y80__R2_CONB_0;
  wire tie_lo_T2Y81__R2_CONB_0;
  wire tie_lo_T2Y82__R2_CONB_0;
  wire tie_lo_T2Y83__R2_CONB_0;
  wire tie_lo_T2Y84__R2_CONB_0;
  wire tie_lo_T2Y85__R2_CONB_0;
  wire tie_lo_T2Y86__R2_CONB_0;
  wire tie_lo_T2Y87__R2_CONB_0;
  wire tie_lo_T2Y88__R2_CONB_0;
  wire tie_lo_T2Y89__R2_CONB_0;
  wire tie_lo_T2Y8__R2_CONB_0;
  wire tie_lo_T2Y9__R2_CONB_0;
  wire tie_lo_T30Y0__R2_CONB_0;
  wire tie_lo_T30Y10__R2_CONB_0;
  wire tie_lo_T30Y11__R2_CONB_0;
  wire tie_lo_T30Y12__R2_CONB_0;
  wire tie_lo_T30Y13__R2_CONB_0;
  wire tie_lo_T30Y14__R2_CONB_0;
  wire tie_lo_T30Y15__R2_CONB_0;
  wire tie_lo_T30Y16__R2_CONB_0;
  wire tie_lo_T30Y17__R2_CONB_0;
  wire tie_lo_T30Y18__R2_CONB_0;
  wire tie_lo_T30Y19__R2_CONB_0;
  wire tie_lo_T30Y1__R2_CONB_0;
  wire tie_lo_T30Y20__R2_CONB_0;
  wire tie_lo_T30Y21__R2_CONB_0;
  wire tie_lo_T30Y22__R2_CONB_0;
  wire tie_lo_T30Y23__R2_CONB_0;
  wire tie_lo_T30Y24__R2_CONB_0;
  wire tie_lo_T30Y25__R2_CONB_0;
  wire tie_lo_T30Y26__R2_CONB_0;
  wire tie_lo_T30Y27__R2_CONB_0;
  wire tie_lo_T30Y28__R2_CONB_0;
  wire tie_lo_T30Y29__R2_CONB_0;
  wire tie_lo_T30Y2__R2_CONB_0;
  wire tie_lo_T30Y30__R2_CONB_0;
  wire tie_lo_T30Y31__R2_CONB_0;
  wire tie_lo_T30Y32__R2_CONB_0;
  wire tie_lo_T30Y33__R2_CONB_0;
  wire tie_lo_T30Y34__R2_CONB_0;
  wire tie_lo_T30Y35__R2_CONB_0;
  wire tie_lo_T30Y36__R2_CONB_0;
  wire tie_lo_T30Y37__R2_CONB_0;
  wire tie_lo_T30Y38__R2_CONB_0;
  wire tie_lo_T30Y39__R2_CONB_0;
  wire tie_lo_T30Y3__R2_CONB_0;
  wire tie_lo_T30Y40__R2_CONB_0;
  wire tie_lo_T30Y41__R2_CONB_0;
  wire tie_lo_T30Y42__R2_CONB_0;
  wire tie_lo_T30Y43__R2_CONB_0;
  wire tie_lo_T30Y44__R2_CONB_0;
  wire tie_lo_T30Y45__R2_CONB_0;
  wire tie_lo_T30Y46__R2_CONB_0;
  wire tie_lo_T30Y47__R2_CONB_0;
  wire tie_lo_T30Y48__R2_CONB_0;
  wire tie_lo_T30Y49__R2_CONB_0;
  wire tie_lo_T30Y4__R2_CONB_0;
  wire tie_lo_T30Y50__R2_CONB_0;
  wire tie_lo_T30Y51__R2_CONB_0;
  wire tie_lo_T30Y52__R2_CONB_0;
  wire tie_lo_T30Y53__R2_CONB_0;
  wire tie_lo_T30Y54__R2_CONB_0;
  wire tie_lo_T30Y55__R2_CONB_0;
  wire tie_lo_T30Y56__R2_CONB_0;
  wire tie_lo_T30Y57__R2_CONB_0;
  wire tie_lo_T30Y58__R2_CONB_0;
  wire tie_lo_T30Y59__R2_CONB_0;
  wire tie_lo_T30Y5__R2_CONB_0;
  wire tie_lo_T30Y60__R2_CONB_0;
  wire tie_lo_T30Y61__R2_CONB_0;
  wire tie_lo_T30Y62__R2_CONB_0;
  wire tie_lo_T30Y63__R2_CONB_0;
  wire tie_lo_T30Y64__R2_CONB_0;
  wire tie_lo_T30Y65__R2_CONB_0;
  wire tie_lo_T30Y66__R2_CONB_0;
  wire tie_lo_T30Y67__R2_CONB_0;
  wire tie_lo_T30Y68__R2_CONB_0;
  wire tie_lo_T30Y69__R2_CONB_0;
  wire tie_lo_T30Y6__R2_CONB_0;
  wire tie_lo_T30Y70__R2_CONB_0;
  wire tie_lo_T30Y71__R2_CONB_0;
  wire tie_lo_T30Y72__R2_CONB_0;
  wire tie_lo_T30Y73__R2_CONB_0;
  wire tie_lo_T30Y74__R2_CONB_0;
  wire tie_lo_T30Y75__R2_CONB_0;
  wire tie_lo_T30Y76__R2_CONB_0;
  wire tie_lo_T30Y77__R2_CONB_0;
  wire tie_lo_T30Y78__R2_CONB_0;
  wire tie_lo_T30Y79__R2_CONB_0;
  wire tie_lo_T30Y7__R2_CONB_0;
  wire tie_lo_T30Y80__R2_CONB_0;
  wire tie_lo_T30Y81__R2_CONB_0;
  wire tie_lo_T30Y82__R2_CONB_0;
  wire tie_lo_T30Y83__R2_CONB_0;
  wire tie_lo_T30Y84__R2_CONB_0;
  wire tie_lo_T30Y85__R2_CONB_0;
  wire tie_lo_T30Y86__R2_CONB_0;
  wire tie_lo_T30Y87__R2_CONB_0;
  wire tie_lo_T30Y88__R2_CONB_0;
  wire tie_lo_T30Y89__R2_CONB_0;
  wire tie_lo_T30Y8__R2_CONB_0;
  wire tie_lo_T30Y9__R2_CONB_0;
  wire tie_lo_T31Y0__R2_CONB_0;
  wire tie_lo_T31Y10__R2_CONB_0;
  wire tie_lo_T31Y11__R2_CONB_0;
  wire tie_lo_T31Y12__R2_CONB_0;
  wire tie_lo_T31Y13__R2_CONB_0;
  wire tie_lo_T31Y14__R2_CONB_0;
  wire tie_lo_T31Y15__R2_CONB_0;
  wire tie_lo_T31Y16__R2_CONB_0;
  wire tie_lo_T31Y17__R2_CONB_0;
  wire tie_lo_T31Y18__R2_CONB_0;
  wire tie_lo_T31Y19__R2_CONB_0;
  wire tie_lo_T31Y1__R2_CONB_0;
  wire tie_lo_T31Y20__R2_CONB_0;
  wire tie_lo_T31Y21__R2_CONB_0;
  wire tie_lo_T31Y22__R2_CONB_0;
  wire tie_lo_T31Y23__R2_CONB_0;
  wire tie_lo_T31Y24__R2_CONB_0;
  wire tie_lo_T31Y25__R2_CONB_0;
  wire tie_lo_T31Y26__R2_CONB_0;
  wire tie_lo_T31Y27__R2_CONB_0;
  wire tie_lo_T31Y28__R2_CONB_0;
  wire tie_lo_T31Y29__R2_CONB_0;
  wire tie_lo_T31Y2__R2_CONB_0;
  wire tie_lo_T31Y30__R2_CONB_0;
  wire tie_lo_T31Y31__R2_CONB_0;
  wire tie_lo_T31Y32__R2_CONB_0;
  wire tie_lo_T31Y33__R2_CONB_0;
  wire tie_lo_T31Y34__R2_CONB_0;
  wire tie_lo_T31Y35__R2_CONB_0;
  wire tie_lo_T31Y36__R2_CONB_0;
  wire tie_lo_T31Y37__R2_CONB_0;
  wire tie_lo_T31Y38__R2_CONB_0;
  wire tie_lo_T31Y39__R2_CONB_0;
  wire tie_lo_T31Y3__R2_CONB_0;
  wire tie_lo_T31Y40__R2_CONB_0;
  wire tie_lo_T31Y41__R2_CONB_0;
  wire tie_lo_T31Y42__R2_CONB_0;
  wire tie_lo_T31Y43__R2_CONB_0;
  wire tie_lo_T31Y44__R2_CONB_0;
  wire tie_lo_T31Y45__R2_CONB_0;
  wire tie_lo_T31Y46__R2_CONB_0;
  wire tie_lo_T31Y47__R2_CONB_0;
  wire tie_lo_T31Y48__R2_CONB_0;
  wire tie_lo_T31Y49__R2_CONB_0;
  wire tie_lo_T31Y4__R2_CONB_0;
  wire tie_lo_T31Y50__R2_CONB_0;
  wire tie_lo_T31Y51__R2_CONB_0;
  wire tie_lo_T31Y52__R2_CONB_0;
  wire tie_lo_T31Y53__R2_CONB_0;
  wire tie_lo_T31Y54__R2_CONB_0;
  wire tie_lo_T31Y55__R2_CONB_0;
  wire tie_lo_T31Y56__R2_CONB_0;
  wire tie_lo_T31Y57__R2_CONB_0;
  wire tie_lo_T31Y58__R2_CONB_0;
  wire tie_lo_T31Y59__R2_CONB_0;
  wire tie_lo_T31Y5__R2_CONB_0;
  wire tie_lo_T31Y60__R2_CONB_0;
  wire tie_lo_T31Y61__R2_CONB_0;
  wire tie_lo_T31Y62__R2_CONB_0;
  wire tie_lo_T31Y63__R2_CONB_0;
  wire tie_lo_T31Y64__R2_CONB_0;
  wire tie_lo_T31Y65__R2_CONB_0;
  wire tie_lo_T31Y66__R2_CONB_0;
  wire tie_lo_T31Y67__R2_CONB_0;
  wire tie_lo_T31Y68__R2_CONB_0;
  wire tie_lo_T31Y69__R2_CONB_0;
  wire tie_lo_T31Y6__R2_CONB_0;
  wire tie_lo_T31Y70__R2_CONB_0;
  wire tie_lo_T31Y71__R2_CONB_0;
  wire tie_lo_T31Y72__R2_CONB_0;
  wire tie_lo_T31Y73__R2_CONB_0;
  wire tie_lo_T31Y74__R2_CONB_0;
  wire tie_lo_T31Y75__R2_CONB_0;
  wire tie_lo_T31Y76__R2_CONB_0;
  wire tie_lo_T31Y77__R2_CONB_0;
  wire tie_lo_T31Y78__R2_CONB_0;
  wire tie_lo_T31Y79__R2_CONB_0;
  wire tie_lo_T31Y7__R2_CONB_0;
  wire tie_lo_T31Y80__R2_CONB_0;
  wire tie_lo_T31Y81__R2_CONB_0;
  wire tie_lo_T31Y82__R2_CONB_0;
  wire tie_lo_T31Y83__R2_CONB_0;
  wire tie_lo_T31Y84__R2_CONB_0;
  wire tie_lo_T31Y85__R2_CONB_0;
  wire tie_lo_T31Y86__R2_CONB_0;
  wire tie_lo_T31Y87__R2_CONB_0;
  wire tie_lo_T31Y88__R2_CONB_0;
  wire tie_lo_T31Y89__R2_CONB_0;
  wire tie_lo_T31Y8__R2_CONB_0;
  wire tie_lo_T31Y9__R2_CONB_0;
  wire tie_lo_T32Y0__R2_CONB_0;
  wire tie_lo_T32Y10__R2_CONB_0;
  wire tie_lo_T32Y11__R2_CONB_0;
  wire tie_lo_T32Y12__R2_CONB_0;
  wire tie_lo_T32Y13__R2_CONB_0;
  wire tie_lo_T32Y14__R2_CONB_0;
  wire tie_lo_T32Y15__R2_CONB_0;
  wire tie_lo_T32Y16__R2_CONB_0;
  wire tie_lo_T32Y17__R2_CONB_0;
  wire tie_lo_T32Y18__R2_CONB_0;
  wire tie_lo_T32Y19__R2_CONB_0;
  wire tie_lo_T32Y1__R2_CONB_0;
  wire tie_lo_T32Y20__R2_CONB_0;
  wire tie_lo_T32Y21__R2_CONB_0;
  wire tie_lo_T32Y22__R2_CONB_0;
  wire tie_lo_T32Y23__R2_CONB_0;
  wire tie_lo_T32Y24__R2_CONB_0;
  wire tie_lo_T32Y25__R2_CONB_0;
  wire tie_lo_T32Y26__R2_CONB_0;
  wire tie_lo_T32Y27__R2_CONB_0;
  wire tie_lo_T32Y28__R2_CONB_0;
  wire tie_lo_T32Y29__R2_CONB_0;
  wire tie_lo_T32Y2__R2_CONB_0;
  wire tie_lo_T32Y30__R2_CONB_0;
  wire tie_lo_T32Y31__R2_CONB_0;
  wire tie_lo_T32Y32__R2_CONB_0;
  wire tie_lo_T32Y33__R2_CONB_0;
  wire tie_lo_T32Y34__R2_CONB_0;
  wire tie_lo_T32Y35__R2_CONB_0;
  wire tie_lo_T32Y36__R2_CONB_0;
  wire tie_lo_T32Y37__R2_CONB_0;
  wire tie_lo_T32Y38__R2_CONB_0;
  wire tie_lo_T32Y39__R2_CONB_0;
  wire tie_lo_T32Y3__R2_CONB_0;
  wire tie_lo_T32Y40__R2_CONB_0;
  wire tie_lo_T32Y41__R2_CONB_0;
  wire tie_lo_T32Y42__R2_CONB_0;
  wire tie_lo_T32Y43__R2_CONB_0;
  wire tie_lo_T32Y44__R2_CONB_0;
  wire tie_lo_T32Y45__R2_CONB_0;
  wire tie_lo_T32Y46__R2_CONB_0;
  wire tie_lo_T32Y47__R2_CONB_0;
  wire tie_lo_T32Y48__R2_CONB_0;
  wire tie_lo_T32Y49__R2_CONB_0;
  wire tie_lo_T32Y4__R2_CONB_0;
  wire tie_lo_T32Y50__R2_CONB_0;
  wire tie_lo_T32Y51__R2_CONB_0;
  wire tie_lo_T32Y52__R2_CONB_0;
  wire tie_lo_T32Y53__R2_CONB_0;
  wire tie_lo_T32Y54__R2_CONB_0;
  wire tie_lo_T32Y55__R2_CONB_0;
  wire tie_lo_T32Y56__R2_CONB_0;
  wire tie_lo_T32Y57__R2_CONB_0;
  wire tie_lo_T32Y58__R2_CONB_0;
  wire tie_lo_T32Y59__R2_CONB_0;
  wire tie_lo_T32Y5__R2_CONB_0;
  wire tie_lo_T32Y60__R2_CONB_0;
  wire tie_lo_T32Y61__R2_CONB_0;
  wire tie_lo_T32Y62__R2_CONB_0;
  wire tie_lo_T32Y63__R2_CONB_0;
  wire tie_lo_T32Y64__R2_CONB_0;
  wire tie_lo_T32Y65__R2_CONB_0;
  wire tie_lo_T32Y66__R2_CONB_0;
  wire tie_lo_T32Y67__R2_CONB_0;
  wire tie_lo_T32Y68__R2_CONB_0;
  wire tie_lo_T32Y69__R2_CONB_0;
  wire tie_lo_T32Y6__R2_CONB_0;
  wire tie_lo_T32Y70__R2_CONB_0;
  wire tie_lo_T32Y71__R2_CONB_0;
  wire tie_lo_T32Y72__R2_CONB_0;
  wire tie_lo_T32Y73__R2_CONB_0;
  wire tie_lo_T32Y74__R2_CONB_0;
  wire tie_lo_T32Y75__R2_CONB_0;
  wire tie_lo_T32Y76__R2_CONB_0;
  wire tie_lo_T32Y77__R2_CONB_0;
  wire tie_lo_T32Y78__R2_CONB_0;
  wire tie_lo_T32Y79__R2_CONB_0;
  wire tie_lo_T32Y7__R2_CONB_0;
  wire tie_lo_T32Y80__R2_CONB_0;
  wire tie_lo_T32Y81__R2_CONB_0;
  wire tie_lo_T32Y82__R2_CONB_0;
  wire tie_lo_T32Y83__R2_CONB_0;
  wire tie_lo_T32Y84__R2_CONB_0;
  wire tie_lo_T32Y85__R2_CONB_0;
  wire tie_lo_T32Y86__R2_CONB_0;
  wire tie_lo_T32Y87__R2_CONB_0;
  wire tie_lo_T32Y88__R2_CONB_0;
  wire tie_lo_T32Y89__R2_CONB_0;
  wire tie_lo_T32Y8__R2_CONB_0;
  wire tie_lo_T32Y9__R2_CONB_0;
  wire tie_lo_T33Y0__R2_CONB_0;
  wire tie_lo_T33Y10__R2_CONB_0;
  wire tie_lo_T33Y11__R2_CONB_0;
  wire tie_lo_T33Y12__R2_CONB_0;
  wire tie_lo_T33Y13__R2_CONB_0;
  wire tie_lo_T33Y14__R2_CONB_0;
  wire tie_lo_T33Y15__R2_CONB_0;
  wire tie_lo_T33Y16__R2_CONB_0;
  wire tie_lo_T33Y17__R2_CONB_0;
  wire tie_lo_T33Y18__R2_CONB_0;
  wire tie_lo_T33Y19__R2_CONB_0;
  wire tie_lo_T33Y1__R2_CONB_0;
  wire tie_lo_T33Y20__R2_CONB_0;
  wire tie_lo_T33Y21__R2_CONB_0;
  wire tie_lo_T33Y22__R2_CONB_0;
  wire tie_lo_T33Y23__R2_CONB_0;
  wire tie_lo_T33Y24__R2_CONB_0;
  wire tie_lo_T33Y25__R2_CONB_0;
  wire tie_lo_T33Y26__R2_CONB_0;
  wire tie_lo_T33Y27__R2_CONB_0;
  wire tie_lo_T33Y28__R2_CONB_0;
  wire tie_lo_T33Y29__R2_CONB_0;
  wire tie_lo_T33Y2__R2_CONB_0;
  wire tie_lo_T33Y30__R2_CONB_0;
  wire tie_lo_T33Y31__R2_CONB_0;
  wire tie_lo_T33Y32__R2_CONB_0;
  wire tie_lo_T33Y33__R2_CONB_0;
  wire tie_lo_T33Y34__R2_CONB_0;
  wire tie_lo_T33Y35__R2_CONB_0;
  wire tie_lo_T33Y36__R2_CONB_0;
  wire tie_lo_T33Y37__R2_CONB_0;
  wire tie_lo_T33Y38__R2_CONB_0;
  wire tie_lo_T33Y39__R2_CONB_0;
  wire tie_lo_T33Y3__R2_CONB_0;
  wire tie_lo_T33Y40__R2_CONB_0;
  wire tie_lo_T33Y41__R2_CONB_0;
  wire tie_lo_T33Y42__R2_CONB_0;
  wire tie_lo_T33Y43__R2_CONB_0;
  wire tie_lo_T33Y44__R2_CONB_0;
  wire tie_lo_T33Y45__R2_CONB_0;
  wire tie_lo_T33Y46__R2_CONB_0;
  wire tie_lo_T33Y47__R2_CONB_0;
  wire tie_lo_T33Y48__R2_CONB_0;
  wire tie_lo_T33Y49__R2_CONB_0;
  wire tie_lo_T33Y4__R2_CONB_0;
  wire tie_lo_T33Y50__R2_CONB_0;
  wire tie_lo_T33Y51__R2_CONB_0;
  wire tie_lo_T33Y52__R2_CONB_0;
  wire tie_lo_T33Y53__R2_CONB_0;
  wire tie_lo_T33Y54__R2_CONB_0;
  wire tie_lo_T33Y55__R2_CONB_0;
  wire tie_lo_T33Y56__R2_CONB_0;
  wire tie_lo_T33Y57__R2_CONB_0;
  wire tie_lo_T33Y58__R2_CONB_0;
  wire tie_lo_T33Y59__R2_CONB_0;
  wire tie_lo_T33Y5__R2_CONB_0;
  wire tie_lo_T33Y60__R2_CONB_0;
  wire tie_lo_T33Y61__R2_CONB_0;
  wire tie_lo_T33Y62__R2_CONB_0;
  wire tie_lo_T33Y63__R2_CONB_0;
  wire tie_lo_T33Y64__R2_CONB_0;
  wire tie_lo_T33Y65__R2_CONB_0;
  wire tie_lo_T33Y66__R2_CONB_0;
  wire tie_lo_T33Y67__R2_CONB_0;
  wire tie_lo_T33Y68__R2_CONB_0;
  wire tie_lo_T33Y69__R2_CONB_0;
  wire tie_lo_T33Y6__R2_CONB_0;
  wire tie_lo_T33Y70__R2_CONB_0;
  wire tie_lo_T33Y71__R2_CONB_0;
  wire tie_lo_T33Y72__R2_CONB_0;
  wire tie_lo_T33Y73__R2_CONB_0;
  wire tie_lo_T33Y74__R2_CONB_0;
  wire tie_lo_T33Y75__R2_CONB_0;
  wire tie_lo_T33Y76__R2_CONB_0;
  wire tie_lo_T33Y77__R2_CONB_0;
  wire tie_lo_T33Y78__R2_CONB_0;
  wire tie_lo_T33Y79__R2_CONB_0;
  wire tie_lo_T33Y7__R2_CONB_0;
  wire tie_lo_T33Y80__R2_CONB_0;
  wire tie_lo_T33Y81__R2_CONB_0;
  wire tie_lo_T33Y82__R2_CONB_0;
  wire tie_lo_T33Y83__R2_CONB_0;
  wire tie_lo_T33Y84__R2_CONB_0;
  wire tie_lo_T33Y85__R2_CONB_0;
  wire tie_lo_T33Y86__R2_CONB_0;
  wire tie_lo_T33Y87__R2_CONB_0;
  wire tie_lo_T33Y88__R2_CONB_0;
  wire tie_lo_T33Y89__R2_CONB_0;
  wire tie_lo_T33Y8__R2_CONB_0;
  wire tie_lo_T33Y9__R2_CONB_0;
  wire tie_lo_T34Y0__R2_CONB_0;
  wire tie_lo_T34Y10__R2_CONB_0;
  wire tie_lo_T34Y11__R2_CONB_0;
  wire tie_lo_T34Y12__R2_CONB_0;
  wire tie_lo_T34Y13__R2_CONB_0;
  wire tie_lo_T34Y14__R2_CONB_0;
  wire tie_lo_T34Y15__R2_CONB_0;
  wire tie_lo_T34Y16__R2_CONB_0;
  wire tie_lo_T34Y17__R2_CONB_0;
  wire tie_lo_T34Y18__R2_CONB_0;
  wire tie_lo_T34Y19__R2_CONB_0;
  wire tie_lo_T34Y1__R2_CONB_0;
  wire tie_lo_T34Y20__R2_CONB_0;
  wire tie_lo_T34Y21__R2_CONB_0;
  wire tie_lo_T34Y22__R2_CONB_0;
  wire tie_lo_T34Y23__R2_CONB_0;
  wire tie_lo_T34Y24__R2_CONB_0;
  wire tie_lo_T34Y25__R2_CONB_0;
  wire tie_lo_T34Y26__R2_CONB_0;
  wire tie_lo_T34Y27__R2_CONB_0;
  wire tie_lo_T34Y28__R2_CONB_0;
  wire tie_lo_T34Y29__R2_CONB_0;
  wire tie_lo_T34Y2__R2_CONB_0;
  wire tie_lo_T34Y30__R2_CONB_0;
  wire tie_lo_T34Y31__R2_CONB_0;
  wire tie_lo_T34Y32__R2_CONB_0;
  wire tie_lo_T34Y33__R2_CONB_0;
  wire tie_lo_T34Y34__R2_CONB_0;
  wire tie_lo_T34Y35__R2_CONB_0;
  wire tie_lo_T34Y36__R2_CONB_0;
  wire tie_lo_T34Y37__R2_CONB_0;
  wire tie_lo_T34Y38__R2_CONB_0;
  wire tie_lo_T34Y39__R2_CONB_0;
  wire tie_lo_T34Y3__R2_CONB_0;
  wire tie_lo_T34Y40__R2_CONB_0;
  wire tie_lo_T34Y41__R2_CONB_0;
  wire tie_lo_T34Y42__R2_CONB_0;
  wire tie_lo_T34Y43__R2_CONB_0;
  wire tie_lo_T34Y44__R2_CONB_0;
  wire tie_lo_T34Y45__R2_CONB_0;
  wire tie_lo_T34Y46__R2_CONB_0;
  wire tie_lo_T34Y47__R2_CONB_0;
  wire tie_lo_T34Y48__R2_CONB_0;
  wire tie_lo_T34Y49__R2_CONB_0;
  wire tie_lo_T34Y4__R2_CONB_0;
  wire tie_lo_T34Y50__R2_CONB_0;
  wire tie_lo_T34Y51__R2_CONB_0;
  wire tie_lo_T34Y52__R2_CONB_0;
  wire tie_lo_T34Y53__R2_CONB_0;
  wire tie_lo_T34Y54__R2_CONB_0;
  wire tie_lo_T34Y55__R2_CONB_0;
  wire tie_lo_T34Y56__R2_CONB_0;
  wire tie_lo_T34Y57__R2_CONB_0;
  wire tie_lo_T34Y58__R2_CONB_0;
  wire tie_lo_T34Y59__R2_CONB_0;
  wire tie_lo_T34Y5__R2_CONB_0;
  wire tie_lo_T34Y60__R2_CONB_0;
  wire tie_lo_T34Y61__R2_CONB_0;
  wire tie_lo_T34Y62__R2_CONB_0;
  wire tie_lo_T34Y63__R2_CONB_0;
  wire tie_lo_T34Y64__R2_CONB_0;
  wire tie_lo_T34Y65__R2_CONB_0;
  wire tie_lo_T34Y66__R2_CONB_0;
  wire tie_lo_T34Y67__R2_CONB_0;
  wire tie_lo_T34Y68__R2_CONB_0;
  wire tie_lo_T34Y69__R2_CONB_0;
  wire tie_lo_T34Y6__R2_CONB_0;
  wire tie_lo_T34Y70__R2_CONB_0;
  wire tie_lo_T34Y71__R2_CONB_0;
  wire tie_lo_T34Y72__R2_CONB_0;
  wire tie_lo_T34Y73__R2_CONB_0;
  wire tie_lo_T34Y74__R2_CONB_0;
  wire tie_lo_T34Y75__R2_CONB_0;
  wire tie_lo_T34Y76__R2_CONB_0;
  wire tie_lo_T34Y77__R2_CONB_0;
  wire tie_lo_T34Y78__R2_CONB_0;
  wire tie_lo_T34Y79__R2_CONB_0;
  wire tie_lo_T34Y7__R2_CONB_0;
  wire tie_lo_T34Y80__R2_CONB_0;
  wire tie_lo_T34Y81__R2_CONB_0;
  wire tie_lo_T34Y82__R2_CONB_0;
  wire tie_lo_T34Y83__R2_CONB_0;
  wire tie_lo_T34Y84__R2_CONB_0;
  wire tie_lo_T34Y85__R2_CONB_0;
  wire tie_lo_T34Y86__R2_CONB_0;
  wire tie_lo_T34Y87__R2_CONB_0;
  wire tie_lo_T34Y88__R2_CONB_0;
  wire tie_lo_T34Y89__R2_CONB_0;
  wire tie_lo_T34Y8__R2_CONB_0;
  wire tie_lo_T34Y9__R2_CONB_0;
  wire tie_lo_T35Y0__R2_CONB_0;
  wire tie_lo_T35Y10__R2_CONB_0;
  wire tie_lo_T35Y11__R2_CONB_0;
  wire tie_lo_T35Y12__R2_CONB_0;
  wire tie_lo_T35Y13__R2_CONB_0;
  wire tie_lo_T35Y14__R2_CONB_0;
  wire tie_lo_T35Y15__R2_CONB_0;
  wire tie_lo_T35Y16__R2_CONB_0;
  wire tie_lo_T35Y17__R2_CONB_0;
  wire tie_lo_T35Y18__R2_CONB_0;
  wire tie_lo_T35Y19__R2_CONB_0;
  wire tie_lo_T35Y1__R2_CONB_0;
  wire tie_lo_T35Y20__R2_CONB_0;
  wire tie_lo_T35Y21__R2_CONB_0;
  wire tie_lo_T35Y22__R2_CONB_0;
  wire tie_lo_T35Y23__R2_CONB_0;
  wire tie_lo_T35Y24__R2_CONB_0;
  wire tie_lo_T35Y25__R2_CONB_0;
  wire tie_lo_T35Y26__R2_CONB_0;
  wire tie_lo_T35Y27__R2_CONB_0;
  wire tie_lo_T35Y28__R2_CONB_0;
  wire tie_lo_T35Y29__R2_CONB_0;
  wire tie_lo_T35Y2__R2_CONB_0;
  wire tie_lo_T35Y30__R2_CONB_0;
  wire tie_lo_T35Y31__R2_CONB_0;
  wire tie_lo_T35Y32__R2_CONB_0;
  wire tie_lo_T35Y33__R2_CONB_0;
  wire tie_lo_T35Y34__R2_CONB_0;
  wire tie_lo_T35Y35__R2_CONB_0;
  wire tie_lo_T35Y36__R2_CONB_0;
  wire tie_lo_T35Y37__R2_CONB_0;
  wire tie_lo_T35Y38__R2_CONB_0;
  wire tie_lo_T35Y39__R2_CONB_0;
  wire tie_lo_T35Y3__R2_CONB_0;
  wire tie_lo_T35Y40__R2_CONB_0;
  wire tie_lo_T35Y41__R2_CONB_0;
  wire tie_lo_T35Y42__R2_CONB_0;
  wire tie_lo_T35Y43__R2_CONB_0;
  wire tie_lo_T35Y44__R2_CONB_0;
  wire tie_lo_T35Y45__R2_CONB_0;
  wire tie_lo_T35Y46__R2_CONB_0;
  wire tie_lo_T35Y47__R2_CONB_0;
  wire tie_lo_T35Y48__R2_CONB_0;
  wire tie_lo_T35Y49__R2_CONB_0;
  wire tie_lo_T35Y4__R2_CONB_0;
  wire tie_lo_T35Y50__R2_CONB_0;
  wire tie_lo_T35Y51__R2_CONB_0;
  wire tie_lo_T35Y52__R2_CONB_0;
  wire tie_lo_T35Y53__R2_CONB_0;
  wire tie_lo_T35Y54__R2_CONB_0;
  wire tie_lo_T35Y55__R2_CONB_0;
  wire tie_lo_T35Y56__R2_CONB_0;
  wire tie_lo_T35Y57__R2_CONB_0;
  wire tie_lo_T35Y58__R2_CONB_0;
  wire tie_lo_T35Y59__R2_CONB_0;
  wire tie_lo_T35Y5__R2_CONB_0;
  wire tie_lo_T35Y60__R2_CONB_0;
  wire tie_lo_T35Y61__R2_CONB_0;
  wire tie_lo_T35Y62__R2_CONB_0;
  wire tie_lo_T35Y63__R2_CONB_0;
  wire tie_lo_T35Y64__R2_CONB_0;
  wire tie_lo_T35Y65__R2_CONB_0;
  wire tie_lo_T35Y66__R2_CONB_0;
  wire tie_lo_T35Y67__R2_CONB_0;
  wire tie_lo_T35Y68__R2_CONB_0;
  wire tie_lo_T35Y69__R2_CONB_0;
  wire tie_lo_T35Y6__R2_CONB_0;
  wire tie_lo_T35Y70__R2_CONB_0;
  wire tie_lo_T35Y71__R2_CONB_0;
  wire tie_lo_T35Y72__R2_CONB_0;
  wire tie_lo_T35Y73__R2_CONB_0;
  wire tie_lo_T35Y74__R2_CONB_0;
  wire tie_lo_T35Y75__R2_CONB_0;
  wire tie_lo_T35Y76__R2_CONB_0;
  wire tie_lo_T35Y77__R2_CONB_0;
  wire tie_lo_T35Y78__R2_CONB_0;
  wire tie_lo_T35Y79__R2_CONB_0;
  wire tie_lo_T35Y7__R2_CONB_0;
  wire tie_lo_T35Y80__R2_CONB_0;
  wire tie_lo_T35Y81__R2_CONB_0;
  wire tie_lo_T35Y82__R2_CONB_0;
  wire tie_lo_T35Y83__R2_CONB_0;
  wire tie_lo_T35Y84__R2_CONB_0;
  wire tie_lo_T35Y85__R2_CONB_0;
  wire tie_lo_T35Y86__R2_CONB_0;
  wire tie_lo_T35Y87__R2_CONB_0;
  wire tie_lo_T35Y88__R2_CONB_0;
  wire tie_lo_T35Y89__R2_CONB_0;
  wire tie_lo_T35Y8__R2_CONB_0;
  wire tie_lo_T35Y9__R2_CONB_0;
  wire tie_lo_T3Y0__R2_CONB_0;
  wire tie_lo_T3Y10__R2_CONB_0;
  wire tie_lo_T3Y11__R2_CONB_0;
  wire tie_lo_T3Y12__R2_CONB_0;
  wire tie_lo_T3Y13__R2_CONB_0;
  wire tie_lo_T3Y14__R2_CONB_0;
  wire tie_lo_T3Y15__R2_CONB_0;
  wire tie_lo_T3Y16__R2_CONB_0;
  wire tie_lo_T3Y17__R2_CONB_0;
  wire tie_lo_T3Y18__R2_CONB_0;
  wire tie_lo_T3Y19__R2_CONB_0;
  wire tie_lo_T3Y1__R2_CONB_0;
  wire tie_lo_T3Y20__R2_CONB_0;
  wire tie_lo_T3Y21__R2_CONB_0;
  wire tie_lo_T3Y22__R2_CONB_0;
  wire tie_lo_T3Y23__R2_CONB_0;
  wire tie_lo_T3Y24__R2_CONB_0;
  wire tie_lo_T3Y25__R2_CONB_0;
  wire tie_lo_T3Y26__R2_CONB_0;
  wire tie_lo_T3Y27__R2_CONB_0;
  wire tie_lo_T3Y28__R2_CONB_0;
  wire tie_lo_T3Y29__R2_CONB_0;
  wire tie_lo_T3Y2__R2_CONB_0;
  wire tie_lo_T3Y30__R2_CONB_0;
  wire tie_lo_T3Y31__R2_CONB_0;
  wire tie_lo_T3Y32__R2_CONB_0;
  wire tie_lo_T3Y33__R2_CONB_0;
  wire tie_lo_T3Y34__R2_CONB_0;
  wire tie_lo_T3Y35__R2_CONB_0;
  wire tie_lo_T3Y36__R2_CONB_0;
  wire tie_lo_T3Y37__R2_CONB_0;
  wire tie_lo_T3Y38__R2_CONB_0;
  wire tie_lo_T3Y39__R2_CONB_0;
  wire tie_lo_T3Y3__R2_CONB_0;
  wire tie_lo_T3Y40__R2_CONB_0;
  wire tie_lo_T3Y41__R2_CONB_0;
  wire tie_lo_T3Y42__R2_CONB_0;
  wire tie_lo_T3Y43__R2_CONB_0;
  wire tie_lo_T3Y44__R2_CONB_0;
  wire tie_lo_T3Y45__R2_CONB_0;
  wire tie_lo_T3Y46__R2_CONB_0;
  wire tie_lo_T3Y47__R2_CONB_0;
  wire tie_lo_T3Y48__R2_CONB_0;
  wire tie_lo_T3Y49__R2_CONB_0;
  wire tie_lo_T3Y4__R2_CONB_0;
  wire tie_lo_T3Y50__R2_CONB_0;
  wire tie_lo_T3Y51__R2_CONB_0;
  wire tie_lo_T3Y52__R2_CONB_0;
  wire tie_lo_T3Y53__R2_CONB_0;
  wire tie_lo_T3Y54__R2_CONB_0;
  wire tie_lo_T3Y55__R2_CONB_0;
  wire tie_lo_T3Y56__R2_CONB_0;
  wire tie_lo_T3Y57__R2_CONB_0;
  wire tie_lo_T3Y58__R2_CONB_0;
  wire tie_lo_T3Y59__R2_CONB_0;
  wire tie_lo_T3Y5__R2_CONB_0;
  wire tie_lo_T3Y60__R2_CONB_0;
  wire tie_lo_T3Y61__R2_CONB_0;
  wire tie_lo_T3Y62__R2_CONB_0;
  wire tie_lo_T3Y63__R2_CONB_0;
  wire tie_lo_T3Y64__R2_CONB_0;
  wire tie_lo_T3Y65__R2_CONB_0;
  wire tie_lo_T3Y66__R2_CONB_0;
  wire tie_lo_T3Y67__R2_CONB_0;
  wire tie_lo_T3Y68__R2_CONB_0;
  wire tie_lo_T3Y69__R2_CONB_0;
  wire tie_lo_T3Y6__R2_CONB_0;
  wire tie_lo_T3Y70__R2_CONB_0;
  wire tie_lo_T3Y71__R2_CONB_0;
  wire tie_lo_T3Y72__R2_CONB_0;
  wire tie_lo_T3Y73__R2_CONB_0;
  wire tie_lo_T3Y74__R2_CONB_0;
  wire tie_lo_T3Y75__R2_CONB_0;
  wire tie_lo_T3Y76__R2_CONB_0;
  wire tie_lo_T3Y77__R2_CONB_0;
  wire tie_lo_T3Y78__R2_CONB_0;
  wire tie_lo_T3Y79__R2_CONB_0;
  wire tie_lo_T3Y7__R2_CONB_0;
  wire tie_lo_T3Y80__R2_CONB_0;
  wire tie_lo_T3Y81__R2_CONB_0;
  wire tie_lo_T3Y82__R2_CONB_0;
  wire tie_lo_T3Y83__R2_CONB_0;
  wire tie_lo_T3Y84__R2_CONB_0;
  wire tie_lo_T3Y85__R2_CONB_0;
  wire tie_lo_T3Y86__R2_CONB_0;
  wire tie_lo_T3Y87__R2_CONB_0;
  wire tie_lo_T3Y88__R2_CONB_0;
  wire tie_lo_T3Y89__R2_CONB_0;
  wire tie_lo_T3Y8__R2_CONB_0;
  wire tie_lo_T3Y9__R2_CONB_0;
  wire tie_lo_T4Y0__R2_CONB_0;
  wire tie_lo_T4Y10__R2_CONB_0;
  wire tie_lo_T4Y11__R2_CONB_0;
  wire tie_lo_T4Y12__R2_CONB_0;
  wire tie_lo_T4Y13__R2_CONB_0;
  wire tie_lo_T4Y14__R2_CONB_0;
  wire tie_lo_T4Y15__R2_CONB_0;
  wire tie_lo_T4Y16__R2_CONB_0;
  wire tie_lo_T4Y17__R2_CONB_0;
  wire tie_lo_T4Y18__R2_CONB_0;
  wire tie_lo_T4Y19__R2_CONB_0;
  wire tie_lo_T4Y1__R2_CONB_0;
  wire tie_lo_T4Y20__R2_CONB_0;
  wire tie_lo_T4Y21__R2_CONB_0;
  wire tie_lo_T4Y22__R2_CONB_0;
  wire tie_lo_T4Y23__R2_CONB_0;
  wire tie_lo_T4Y24__R2_CONB_0;
  wire tie_lo_T4Y25__R2_CONB_0;
  wire tie_lo_T4Y26__R2_CONB_0;
  wire tie_lo_T4Y27__R2_CONB_0;
  wire tie_lo_T4Y28__R2_CONB_0;
  wire tie_lo_T4Y29__R2_CONB_0;
  wire tie_lo_T4Y2__R2_CONB_0;
  wire tie_lo_T4Y30__R2_CONB_0;
  wire tie_lo_T4Y31__R2_CONB_0;
  wire tie_lo_T4Y32__R2_CONB_0;
  wire tie_lo_T4Y33__R2_CONB_0;
  wire tie_lo_T4Y34__R2_CONB_0;
  wire tie_lo_T4Y35__R2_CONB_0;
  wire tie_lo_T4Y36__R2_CONB_0;
  wire tie_lo_T4Y37__R2_CONB_0;
  wire tie_lo_T4Y38__R2_CONB_0;
  wire tie_lo_T4Y39__R2_CONB_0;
  wire tie_lo_T4Y3__R2_CONB_0;
  wire tie_lo_T4Y40__R2_CONB_0;
  wire tie_lo_T4Y41__R2_CONB_0;
  wire tie_lo_T4Y42__R2_CONB_0;
  wire tie_lo_T4Y43__R2_CONB_0;
  wire tie_lo_T4Y44__R2_CONB_0;
  wire tie_lo_T4Y45__R2_CONB_0;
  wire tie_lo_T4Y46__R2_CONB_0;
  wire tie_lo_T4Y47__R2_CONB_0;
  wire tie_lo_T4Y48__R2_CONB_0;
  wire tie_lo_T4Y49__R2_CONB_0;
  wire tie_lo_T4Y4__R2_CONB_0;
  wire tie_lo_T4Y50__R2_CONB_0;
  wire tie_lo_T4Y51__R2_CONB_0;
  wire tie_lo_T4Y52__R2_CONB_0;
  wire tie_lo_T4Y53__R2_CONB_0;
  wire tie_lo_T4Y54__R2_CONB_0;
  wire tie_lo_T4Y55__R2_CONB_0;
  wire tie_lo_T4Y56__R2_CONB_0;
  wire tie_lo_T4Y57__R2_CONB_0;
  wire tie_lo_T4Y58__R2_CONB_0;
  wire tie_lo_T4Y59__R2_CONB_0;
  wire tie_lo_T4Y5__R2_CONB_0;
  wire tie_lo_T4Y60__R2_CONB_0;
  wire tie_lo_T4Y61__R2_CONB_0;
  wire tie_lo_T4Y62__R2_CONB_0;
  wire tie_lo_T4Y63__R2_CONB_0;
  wire tie_lo_T4Y64__R2_CONB_0;
  wire tie_lo_T4Y65__R2_CONB_0;
  wire tie_lo_T4Y66__R2_CONB_0;
  wire tie_lo_T4Y67__R2_CONB_0;
  wire tie_lo_T4Y68__R2_CONB_0;
  wire tie_lo_T4Y69__R2_CONB_0;
  wire tie_lo_T4Y6__R2_CONB_0;
  wire tie_lo_T4Y70__R2_CONB_0;
  wire tie_lo_T4Y71__R2_CONB_0;
  wire tie_lo_T4Y72__R2_CONB_0;
  wire tie_lo_T4Y73__R2_CONB_0;
  wire tie_lo_T4Y74__R2_CONB_0;
  wire tie_lo_T4Y75__R2_CONB_0;
  wire tie_lo_T4Y76__R2_CONB_0;
  wire tie_lo_T4Y77__R2_CONB_0;
  wire tie_lo_T4Y78__R2_CONB_0;
  wire tie_lo_T4Y79__R2_CONB_0;
  wire tie_lo_T4Y7__R2_CONB_0;
  wire tie_lo_T4Y80__R2_CONB_0;
  wire tie_lo_T4Y81__R2_CONB_0;
  wire tie_lo_T4Y82__R2_CONB_0;
  wire tie_lo_T4Y83__R2_CONB_0;
  wire tie_lo_T4Y84__R2_CONB_0;
  wire tie_lo_T4Y85__R2_CONB_0;
  wire tie_lo_T4Y86__R2_CONB_0;
  wire tie_lo_T4Y87__R2_CONB_0;
  wire tie_lo_T4Y88__R2_CONB_0;
  wire tie_lo_T4Y89__R2_CONB_0;
  wire tie_lo_T4Y8__R2_CONB_0;
  wire tie_lo_T4Y9__R2_CONB_0;
  wire tie_lo_T5Y0__R2_CONB_0;
  wire tie_lo_T5Y10__R2_CONB_0;
  wire tie_lo_T5Y11__R2_CONB_0;
  wire tie_lo_T5Y12__R2_CONB_0;
  wire tie_lo_T5Y13__R2_CONB_0;
  wire tie_lo_T5Y14__R2_CONB_0;
  wire tie_lo_T5Y15__R2_CONB_0;
  wire tie_lo_T5Y16__R2_CONB_0;
  wire tie_lo_T5Y17__R2_CONB_0;
  wire tie_lo_T5Y18__R2_CONB_0;
  wire tie_lo_T5Y19__R2_CONB_0;
  wire tie_lo_T5Y1__R2_CONB_0;
  wire tie_lo_T5Y20__R2_CONB_0;
  wire tie_lo_T5Y21__R2_CONB_0;
  wire tie_lo_T5Y22__R2_CONB_0;
  wire tie_lo_T5Y23__R2_CONB_0;
  wire tie_lo_T5Y24__R2_CONB_0;
  wire tie_lo_T5Y25__R2_CONB_0;
  wire tie_lo_T5Y26__R2_CONB_0;
  wire tie_lo_T5Y27__R2_CONB_0;
  wire tie_lo_T5Y28__R2_CONB_0;
  wire tie_lo_T5Y29__R2_CONB_0;
  wire tie_lo_T5Y2__R2_CONB_0;
  wire tie_lo_T5Y30__R2_CONB_0;
  wire tie_lo_T5Y31__R2_CONB_0;
  wire tie_lo_T5Y32__R2_CONB_0;
  wire tie_lo_T5Y33__R2_CONB_0;
  wire tie_lo_T5Y34__R2_CONB_0;
  wire tie_lo_T5Y35__R2_CONB_0;
  wire tie_lo_T5Y36__R2_CONB_0;
  wire tie_lo_T5Y37__R2_CONB_0;
  wire tie_lo_T5Y38__R2_CONB_0;
  wire tie_lo_T5Y39__R2_CONB_0;
  wire tie_lo_T5Y3__R2_CONB_0;
  wire tie_lo_T5Y40__R2_CONB_0;
  wire tie_lo_T5Y41__R2_CONB_0;
  wire tie_lo_T5Y42__R2_CONB_0;
  wire tie_lo_T5Y43__R2_CONB_0;
  wire tie_lo_T5Y44__R2_CONB_0;
  wire tie_lo_T5Y45__R2_CONB_0;
  wire tie_lo_T5Y46__R2_CONB_0;
  wire tie_lo_T5Y47__R2_CONB_0;
  wire tie_lo_T5Y48__R2_CONB_0;
  wire tie_lo_T5Y49__R2_CONB_0;
  wire tie_lo_T5Y4__R2_CONB_0;
  wire tie_lo_T5Y50__R2_CONB_0;
  wire tie_lo_T5Y51__R2_CONB_0;
  wire tie_lo_T5Y52__R2_CONB_0;
  wire tie_lo_T5Y53__R2_CONB_0;
  wire tie_lo_T5Y54__R2_CONB_0;
  wire tie_lo_T5Y55__R2_CONB_0;
  wire tie_lo_T5Y56__R2_CONB_0;
  wire tie_lo_T5Y57__R2_CONB_0;
  wire tie_lo_T5Y58__R2_CONB_0;
  wire tie_lo_T5Y59__R2_CONB_0;
  wire tie_lo_T5Y5__R2_CONB_0;
  wire tie_lo_T5Y60__R2_CONB_0;
  wire tie_lo_T5Y61__R2_CONB_0;
  wire tie_lo_T5Y62__R2_CONB_0;
  wire tie_lo_T5Y63__R2_CONB_0;
  wire tie_lo_T5Y64__R2_CONB_0;
  wire tie_lo_T5Y65__R2_CONB_0;
  wire tie_lo_T5Y66__R2_CONB_0;
  wire tie_lo_T5Y67__R2_CONB_0;
  wire tie_lo_T5Y68__R2_CONB_0;
  wire tie_lo_T5Y69__R2_CONB_0;
  wire tie_lo_T5Y6__R2_CONB_0;
  wire tie_lo_T5Y70__R2_CONB_0;
  wire tie_lo_T5Y71__R2_CONB_0;
  wire tie_lo_T5Y72__R2_CONB_0;
  wire tie_lo_T5Y73__R2_CONB_0;
  wire tie_lo_T5Y74__R2_CONB_0;
  wire tie_lo_T5Y75__R2_CONB_0;
  wire tie_lo_T5Y76__R2_CONB_0;
  wire tie_lo_T5Y77__R2_CONB_0;
  wire tie_lo_T5Y78__R2_CONB_0;
  wire tie_lo_T5Y79__R2_CONB_0;
  wire tie_lo_T5Y7__R2_CONB_0;
  wire tie_lo_T5Y80__R2_CONB_0;
  wire tie_lo_T5Y81__R2_CONB_0;
  wire tie_lo_T5Y82__R2_CONB_0;
  wire tie_lo_T5Y83__R2_CONB_0;
  wire tie_lo_T5Y84__R2_CONB_0;
  wire tie_lo_T5Y85__R2_CONB_0;
  wire tie_lo_T5Y86__R2_CONB_0;
  wire tie_lo_T5Y87__R2_CONB_0;
  wire tie_lo_T5Y88__R2_CONB_0;
  wire tie_lo_T5Y89__R2_CONB_0;
  wire tie_lo_T5Y8__R2_CONB_0;
  wire tie_lo_T5Y9__R2_CONB_0;
  wire tie_lo_T6Y0__R2_CONB_0;
  wire tie_lo_T6Y10__R2_CONB_0;
  wire tie_lo_T6Y11__R2_CONB_0;
  wire tie_lo_T6Y12__R2_CONB_0;
  wire tie_lo_T6Y13__R2_CONB_0;
  wire tie_lo_T6Y14__R2_CONB_0;
  wire tie_lo_T6Y15__R2_CONB_0;
  wire tie_lo_T6Y16__R2_CONB_0;
  wire tie_lo_T6Y17__R2_CONB_0;
  wire tie_lo_T6Y18__R2_CONB_0;
  wire tie_lo_T6Y19__R2_CONB_0;
  wire tie_lo_T6Y1__R2_CONB_0;
  wire tie_lo_T6Y20__R2_CONB_0;
  wire tie_lo_T6Y21__R2_CONB_0;
  wire tie_lo_T6Y22__R2_CONB_0;
  wire tie_lo_T6Y23__R2_CONB_0;
  wire tie_lo_T6Y24__R2_CONB_0;
  wire tie_lo_T6Y25__R2_CONB_0;
  wire tie_lo_T6Y26__R2_CONB_0;
  wire tie_lo_T6Y27__R2_CONB_0;
  wire tie_lo_T6Y28__R2_CONB_0;
  wire tie_lo_T6Y29__R2_CONB_0;
  wire tie_lo_T6Y2__R2_CONB_0;
  wire tie_lo_T6Y30__R2_CONB_0;
  wire tie_lo_T6Y31__R2_CONB_0;
  wire tie_lo_T6Y32__R2_CONB_0;
  wire tie_lo_T6Y33__R2_CONB_0;
  wire tie_lo_T6Y34__R2_CONB_0;
  wire tie_lo_T6Y35__R2_CONB_0;
  wire tie_lo_T6Y36__R2_CONB_0;
  wire tie_lo_T6Y37__R2_CONB_0;
  wire tie_lo_T6Y38__R2_CONB_0;
  wire tie_lo_T6Y39__R2_CONB_0;
  wire tie_lo_T6Y3__R2_CONB_0;
  wire tie_lo_T6Y40__R2_CONB_0;
  wire tie_lo_T6Y41__R2_CONB_0;
  wire tie_lo_T6Y42__R2_CONB_0;
  wire tie_lo_T6Y43__R2_CONB_0;
  wire tie_lo_T6Y44__R2_CONB_0;
  wire tie_lo_T6Y45__R2_CONB_0;
  wire tie_lo_T6Y46__R2_CONB_0;
  wire tie_lo_T6Y47__R2_CONB_0;
  wire tie_lo_T6Y48__R2_CONB_0;
  wire tie_lo_T6Y49__R2_CONB_0;
  wire tie_lo_T6Y4__R2_CONB_0;
  wire tie_lo_T6Y50__R2_CONB_0;
  wire tie_lo_T6Y51__R2_CONB_0;
  wire tie_lo_T6Y52__R2_CONB_0;
  wire tie_lo_T6Y53__R2_CONB_0;
  wire tie_lo_T6Y54__R2_CONB_0;
  wire tie_lo_T6Y55__R2_CONB_0;
  wire tie_lo_T6Y56__R2_CONB_0;
  wire tie_lo_T6Y57__R2_CONB_0;
  wire tie_lo_T6Y58__R2_CONB_0;
  wire tie_lo_T6Y59__R2_CONB_0;
  wire tie_lo_T6Y5__R2_CONB_0;
  wire tie_lo_T6Y60__R2_CONB_0;
  wire tie_lo_T6Y61__R2_CONB_0;
  wire tie_lo_T6Y62__R2_CONB_0;
  wire tie_lo_T6Y63__R2_CONB_0;
  wire tie_lo_T6Y64__R2_CONB_0;
  wire tie_lo_T6Y65__R2_CONB_0;
  wire tie_lo_T6Y66__R2_CONB_0;
  wire tie_lo_T6Y67__R2_CONB_0;
  wire tie_lo_T6Y68__R2_CONB_0;
  wire tie_lo_T6Y69__R2_CONB_0;
  wire tie_lo_T6Y6__R2_CONB_0;
  wire tie_lo_T6Y70__R2_CONB_0;
  wire tie_lo_T6Y71__R2_CONB_0;
  wire tie_lo_T6Y72__R2_CONB_0;
  wire tie_lo_T6Y73__R2_CONB_0;
  wire tie_lo_T6Y74__R2_CONB_0;
  wire tie_lo_T6Y75__R2_CONB_0;
  wire tie_lo_T6Y76__R2_CONB_0;
  wire tie_lo_T6Y77__R2_CONB_0;
  wire tie_lo_T6Y78__R2_CONB_0;
  wire tie_lo_T6Y79__R2_CONB_0;
  wire tie_lo_T6Y7__R2_CONB_0;
  wire tie_lo_T6Y80__R2_CONB_0;
  wire tie_lo_T6Y81__R2_CONB_0;
  wire tie_lo_T6Y82__R2_CONB_0;
  wire tie_lo_T6Y83__R2_CONB_0;
  wire tie_lo_T6Y84__R2_CONB_0;
  wire tie_lo_T6Y85__R2_CONB_0;
  wire tie_lo_T6Y86__R2_CONB_0;
  wire tie_lo_T6Y87__R2_CONB_0;
  wire tie_lo_T6Y88__R2_CONB_0;
  wire tie_lo_T6Y89__R2_CONB_0;
  wire tie_lo_T6Y8__R2_CONB_0;
  wire tie_lo_T6Y9__R2_CONB_0;
  wire tie_lo_T7Y0__R2_CONB_0;
  wire tie_lo_T7Y10__R2_CONB_0;
  wire tie_lo_T7Y11__R2_CONB_0;
  wire tie_lo_T7Y12__R2_CONB_0;
  wire tie_lo_T7Y13__R2_CONB_0;
  wire tie_lo_T7Y14__R2_CONB_0;
  wire tie_lo_T7Y15__R2_CONB_0;
  wire tie_lo_T7Y16__R2_CONB_0;
  wire tie_lo_T7Y17__R2_CONB_0;
  wire tie_lo_T7Y18__R2_CONB_0;
  wire tie_lo_T7Y19__R2_CONB_0;
  wire tie_lo_T7Y1__R2_CONB_0;
  wire tie_lo_T7Y20__R2_CONB_0;
  wire tie_lo_T7Y21__R2_CONB_0;
  wire tie_lo_T7Y22__R2_CONB_0;
  wire tie_lo_T7Y23__R2_CONB_0;
  wire tie_lo_T7Y24__R2_CONB_0;
  wire tie_lo_T7Y25__R2_CONB_0;
  wire tie_lo_T7Y26__R2_CONB_0;
  wire tie_lo_T7Y27__R2_CONB_0;
  wire tie_lo_T7Y28__R2_CONB_0;
  wire tie_lo_T7Y29__R2_CONB_0;
  wire tie_lo_T7Y2__R2_CONB_0;
  wire tie_lo_T7Y30__R2_CONB_0;
  wire tie_lo_T7Y31__R2_CONB_0;
  wire tie_lo_T7Y32__R2_CONB_0;
  wire tie_lo_T7Y33__R2_CONB_0;
  wire tie_lo_T7Y34__R2_CONB_0;
  wire tie_lo_T7Y35__R2_CONB_0;
  wire tie_lo_T7Y36__R2_CONB_0;
  wire tie_lo_T7Y37__R2_CONB_0;
  wire tie_lo_T7Y38__R2_CONB_0;
  wire tie_lo_T7Y39__R2_CONB_0;
  wire tie_lo_T7Y3__R2_CONB_0;
  wire tie_lo_T7Y40__R2_CONB_0;
  wire tie_lo_T7Y41__R2_CONB_0;
  wire tie_lo_T7Y42__R2_CONB_0;
  wire tie_lo_T7Y43__R2_CONB_0;
  wire tie_lo_T7Y44__R2_CONB_0;
  wire tie_lo_T7Y45__R2_CONB_0;
  wire tie_lo_T7Y46__R2_CONB_0;
  wire tie_lo_T7Y47__R2_CONB_0;
  wire tie_lo_T7Y48__R2_CONB_0;
  wire tie_lo_T7Y49__R2_CONB_0;
  wire tie_lo_T7Y4__R2_CONB_0;
  wire tie_lo_T7Y50__R2_CONB_0;
  wire tie_lo_T7Y51__R2_CONB_0;
  wire tie_lo_T7Y52__R2_CONB_0;
  wire tie_lo_T7Y53__R2_CONB_0;
  wire tie_lo_T7Y54__R2_CONB_0;
  wire tie_lo_T7Y55__R2_CONB_0;
  wire tie_lo_T7Y56__R2_CONB_0;
  wire tie_lo_T7Y57__R2_CONB_0;
  wire tie_lo_T7Y58__R2_CONB_0;
  wire tie_lo_T7Y59__R2_CONB_0;
  wire tie_lo_T7Y5__R2_CONB_0;
  wire tie_lo_T7Y60__R2_CONB_0;
  wire tie_lo_T7Y61__R2_CONB_0;
  wire tie_lo_T7Y62__R2_CONB_0;
  wire tie_lo_T7Y63__R2_CONB_0;
  wire tie_lo_T7Y64__R2_CONB_0;
  wire tie_lo_T7Y65__R2_CONB_0;
  wire tie_lo_T7Y66__R2_CONB_0;
  wire tie_lo_T7Y67__R2_CONB_0;
  wire tie_lo_T7Y68__R2_CONB_0;
  wire tie_lo_T7Y69__R2_CONB_0;
  wire tie_lo_T7Y6__R2_CONB_0;
  wire tie_lo_T7Y70__R2_CONB_0;
  wire tie_lo_T7Y71__R2_CONB_0;
  wire tie_lo_T7Y72__R2_CONB_0;
  wire tie_lo_T7Y73__R2_CONB_0;
  wire tie_lo_T7Y74__R2_CONB_0;
  wire tie_lo_T7Y75__R2_CONB_0;
  wire tie_lo_T7Y76__R2_CONB_0;
  wire tie_lo_T7Y77__R2_CONB_0;
  wire tie_lo_T7Y78__R2_CONB_0;
  wire tie_lo_T7Y79__R2_CONB_0;
  wire tie_lo_T7Y7__R2_CONB_0;
  wire tie_lo_T7Y80__R2_CONB_0;
  wire tie_lo_T7Y81__R2_CONB_0;
  wire tie_lo_T7Y82__R2_CONB_0;
  wire tie_lo_T7Y83__R2_CONB_0;
  wire tie_lo_T7Y84__R2_CONB_0;
  wire tie_lo_T7Y85__R2_CONB_0;
  wire tie_lo_T7Y86__R2_CONB_0;
  wire tie_lo_T7Y87__R2_CONB_0;
  wire tie_lo_T7Y88__R2_CONB_0;
  wire tie_lo_T7Y89__R2_CONB_0;
  wire tie_lo_T7Y8__R2_CONB_0;
  wire tie_lo_T7Y9__R2_CONB_0;
  wire tie_lo_T8Y0__R2_CONB_0;
  wire tie_lo_T8Y10__R2_CONB_0;
  wire tie_lo_T8Y11__R2_CONB_0;
  wire tie_lo_T8Y12__R2_CONB_0;
  wire tie_lo_T8Y13__R2_CONB_0;
  wire tie_lo_T8Y14__R2_CONB_0;
  wire tie_lo_T8Y15__R2_CONB_0;
  wire tie_lo_T8Y16__R2_CONB_0;
  wire tie_lo_T8Y17__R2_CONB_0;
  wire tie_lo_T8Y18__R2_CONB_0;
  wire tie_lo_T8Y19__R2_CONB_0;
  wire tie_lo_T8Y1__R2_CONB_0;
  wire tie_lo_T8Y20__R2_CONB_0;
  wire tie_lo_T8Y21__R2_CONB_0;
  wire tie_lo_T8Y22__R2_CONB_0;
  wire tie_lo_T8Y23__R2_CONB_0;
  wire tie_lo_T8Y24__R2_CONB_0;
  wire tie_lo_T8Y25__R2_CONB_0;
  wire tie_lo_T8Y26__R2_CONB_0;
  wire tie_lo_T8Y27__R2_CONB_0;
  wire tie_lo_T8Y28__R2_CONB_0;
  wire tie_lo_T8Y29__R2_CONB_0;
  wire tie_lo_T8Y2__R2_CONB_0;
  wire tie_lo_T8Y30__R2_CONB_0;
  wire tie_lo_T8Y31__R2_CONB_0;
  wire tie_lo_T8Y32__R2_CONB_0;
  wire tie_lo_T8Y33__R2_CONB_0;
  wire tie_lo_T8Y34__R2_CONB_0;
  wire tie_lo_T8Y35__R2_CONB_0;
  wire tie_lo_T8Y36__R2_CONB_0;
  wire tie_lo_T8Y37__R2_CONB_0;
  wire tie_lo_T8Y38__R2_CONB_0;
  wire tie_lo_T8Y39__R2_CONB_0;
  wire tie_lo_T8Y3__R2_CONB_0;
  wire tie_lo_T8Y40__R2_CONB_0;
  wire tie_lo_T8Y41__R2_CONB_0;
  wire tie_lo_T8Y42__R2_CONB_0;
  wire tie_lo_T8Y43__R2_CONB_0;
  wire tie_lo_T8Y44__R2_CONB_0;
  wire tie_lo_T8Y45__R2_CONB_0;
  wire tie_lo_T8Y46__R2_CONB_0;
  wire tie_lo_T8Y47__R2_CONB_0;
  wire tie_lo_T8Y48__R2_CONB_0;
  wire tie_lo_T8Y49__R2_CONB_0;
  wire tie_lo_T8Y4__R2_CONB_0;
  wire tie_lo_T8Y50__R2_CONB_0;
  wire tie_lo_T8Y51__R2_CONB_0;
  wire tie_lo_T8Y52__R2_CONB_0;
  wire tie_lo_T8Y53__R2_CONB_0;
  wire tie_lo_T8Y54__R2_CONB_0;
  wire tie_lo_T8Y55__R2_CONB_0;
  wire tie_lo_T8Y56__R2_CONB_0;
  wire tie_lo_T8Y57__R2_CONB_0;
  wire tie_lo_T8Y58__R2_CONB_0;
  wire tie_lo_T8Y59__R2_CONB_0;
  wire tie_lo_T8Y5__R2_CONB_0;
  wire tie_lo_T8Y60__R2_CONB_0;
  wire tie_lo_T8Y61__R2_CONB_0;
  wire tie_lo_T8Y62__R2_CONB_0;
  wire tie_lo_T8Y63__R2_CONB_0;
  wire tie_lo_T8Y64__R2_CONB_0;
  wire tie_lo_T8Y65__R2_CONB_0;
  wire tie_lo_T8Y66__R2_CONB_0;
  wire tie_lo_T8Y67__R2_CONB_0;
  wire tie_lo_T8Y68__R2_CONB_0;
  wire tie_lo_T8Y69__R2_CONB_0;
  wire tie_lo_T8Y6__R2_CONB_0;
  wire tie_lo_T8Y70__R2_CONB_0;
  wire tie_lo_T8Y71__R2_CONB_0;
  wire tie_lo_T8Y72__R2_CONB_0;
  wire tie_lo_T8Y73__R2_CONB_0;
  wire tie_lo_T8Y74__R2_CONB_0;
  wire tie_lo_T8Y75__R2_CONB_0;
  wire tie_lo_T8Y76__R2_CONB_0;
  wire tie_lo_T8Y77__R2_CONB_0;
  wire tie_lo_T8Y78__R2_CONB_0;
  wire tie_lo_T8Y79__R2_CONB_0;
  wire tie_lo_T8Y7__R2_CONB_0;
  wire tie_lo_T8Y80__R2_CONB_0;
  wire tie_lo_T8Y81__R2_CONB_0;
  wire tie_lo_T8Y82__R2_CONB_0;
  wire tie_lo_T8Y83__R2_CONB_0;
  wire tie_lo_T8Y84__R2_CONB_0;
  wire tie_lo_T8Y85__R2_CONB_0;
  wire tie_lo_T8Y86__R2_CONB_0;
  wire tie_lo_T8Y87__R2_CONB_0;
  wire tie_lo_T8Y88__R2_CONB_0;
  wire tie_lo_T8Y89__R2_CONB_0;
  wire tie_lo_T8Y8__R2_CONB_0;
  wire tie_lo_T8Y9__R2_CONB_0;
  wire tie_lo_T9Y0__R2_CONB_0;
  wire tie_lo_T9Y10__R2_CONB_0;
  wire tie_lo_T9Y11__R2_CONB_0;
  wire tie_lo_T9Y12__R2_CONB_0;
  wire tie_lo_T9Y13__R2_CONB_0;
  wire tie_lo_T9Y14__R2_CONB_0;
  wire tie_lo_T9Y15__R2_CONB_0;
  wire tie_lo_T9Y16__R2_CONB_0;
  wire tie_lo_T9Y17__R2_CONB_0;
  wire tie_lo_T9Y18__R2_CONB_0;
  wire tie_lo_T9Y19__R2_CONB_0;
  wire tie_lo_T9Y1__R2_CONB_0;
  wire tie_lo_T9Y20__R2_CONB_0;
  wire tie_lo_T9Y21__R2_CONB_0;
  wire tie_lo_T9Y22__R2_CONB_0;
  wire tie_lo_T9Y23__R2_CONB_0;
  wire tie_lo_T9Y24__R2_CONB_0;
  wire tie_lo_T9Y25__R2_CONB_0;
  wire tie_lo_T9Y26__R2_CONB_0;
  wire tie_lo_T9Y27__R2_CONB_0;
  wire tie_lo_T9Y28__R2_CONB_0;
  wire tie_lo_T9Y29__R2_CONB_0;
  wire tie_lo_T9Y2__R2_CONB_0;
  wire tie_lo_T9Y30__R2_CONB_0;
  wire tie_lo_T9Y31__R2_CONB_0;
  wire tie_lo_T9Y32__R2_CONB_0;
  wire tie_lo_T9Y33__R2_CONB_0;
  wire tie_lo_T9Y34__R2_CONB_0;
  wire tie_lo_T9Y35__R2_CONB_0;
  wire tie_lo_T9Y36__R2_CONB_0;
  wire tie_lo_T9Y37__R2_CONB_0;
  wire tie_lo_T9Y38__R2_CONB_0;
  wire tie_lo_T9Y39__R2_CONB_0;
  wire tie_lo_T9Y3__R2_CONB_0;
  wire tie_lo_T9Y40__R2_CONB_0;
  wire tie_lo_T9Y41__R2_CONB_0;
  wire tie_lo_T9Y42__R2_CONB_0;
  wire tie_lo_T9Y43__R2_CONB_0;
  wire tie_lo_T9Y44__R2_CONB_0;
  wire tie_lo_T9Y45__R2_CONB_0;
  wire tie_lo_T9Y46__R2_CONB_0;
  wire tie_lo_T9Y47__R2_CONB_0;
  wire tie_lo_T9Y48__R2_CONB_0;
  wire tie_lo_T9Y49__R2_CONB_0;
  wire tie_lo_T9Y4__R2_CONB_0;
  wire tie_lo_T9Y50__R2_CONB_0;
  wire tie_lo_T9Y51__R2_CONB_0;
  wire tie_lo_T9Y52__R2_CONB_0;
  wire tie_lo_T9Y53__R2_CONB_0;
  wire tie_lo_T9Y54__R2_CONB_0;
  wire tie_lo_T9Y55__R2_CONB_0;
  wire tie_lo_T9Y56__R2_CONB_0;
  wire tie_lo_T9Y57__R2_CONB_0;
  wire tie_lo_T9Y58__R2_CONB_0;
  wire tie_lo_T9Y59__R2_CONB_0;
  wire tie_lo_T9Y5__R2_CONB_0;
  wire tie_lo_T9Y60__R2_CONB_0;
  wire tie_lo_T9Y61__R2_CONB_0;
  wire tie_lo_T9Y62__R2_CONB_0;
  wire tie_lo_T9Y63__R2_CONB_0;
  wire tie_lo_T9Y64__R2_CONB_0;
  wire tie_lo_T9Y65__R2_CONB_0;
  wire tie_lo_T9Y66__R2_CONB_0;
  wire tie_lo_T9Y67__R2_CONB_0;
  wire tie_lo_T9Y68__R2_CONB_0;
  wire tie_lo_T9Y69__R2_CONB_0;
  wire tie_lo_T9Y6__R2_CONB_0;
  wire tie_lo_T9Y70__R2_CONB_0;
  wire tie_lo_T9Y71__R2_CONB_0;
  wire tie_lo_T9Y72__R2_CONB_0;
  wire tie_lo_T9Y73__R2_CONB_0;
  wire tie_lo_T9Y74__R2_CONB_0;
  wire tie_lo_T9Y75__R2_CONB_0;
  wire tie_lo_T9Y76__R2_CONB_0;
  wire tie_lo_T9Y77__R2_CONB_0;
  wire tie_lo_T9Y78__R2_CONB_0;
  wire tie_lo_T9Y79__R2_CONB_0;
  wire tie_lo_T9Y7__R2_CONB_0;
  wire tie_lo_T9Y80__R2_CONB_0;
  wire tie_lo_T9Y81__R2_CONB_0;
  wire tie_lo_T9Y82__R2_CONB_0;
  wire tie_lo_T9Y83__R2_CONB_0;
  wire tie_lo_T9Y84__R2_CONB_0;
  wire tie_lo_T9Y85__R2_CONB_0;
  wire tie_lo_T9Y86__R2_CONB_0;
  wire tie_lo_T9Y87__R2_CONB_0;
  wire tie_lo_T9Y88__R2_CONB_0;
  wire tie_lo_T9Y89__R2_CONB_0;
  wire tie_lo_T9Y8__R2_CONB_0;
  wire tie_lo_T9Y9__R2_CONB_0;

  // Cell instantiations
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10000 (.A([124]), .B([125]), .X([126]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10001 (.A([127]), .B([126]), .X([128]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10002 (.A([128]), .Y([129]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10003 (.A([130]), .B([129]), .Y([131]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10004 (.A([132]), .B([131]), .Y([133]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10005 (.A([133]), .Y([134]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10006 (.A([132]), .B([131]), .X([135]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10007 (.A([133]), .B([135]), .Y([136]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10008 (.A([39]), .B([136]), .Y([137]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10009 (.A([39]), .B([138]), .X([139]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10010 (.A([137]), .B([139]), .Y([140]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10011 (.A([140]), .Y([141]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10012 (.A([142]), .B([143]), .Y([144]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10013 (.A([145]), .B([146]), .Y([147]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10014 (.A([145]), .B([148]), .Y([149]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10015 (.A([150]), .B([149]), .Y([151]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10016 (.A([152]), .B([153]), .Y([154]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10017 (.A([147]), .B([154]), .Y([155]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10018 (.A([151]), .B([155]), .X([156]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10019 (.A([156]), .Y([157]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10020 (.A([144]), .B([157]), .Y([158]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10021 (.A([134]), .B([158]), .Y([159]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10022 (.A([159]), .Y([160]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10023 (.A([134]), .B([158]), .X([161]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10024 (.A([159]), .B([161]), .Y([162]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10025 (.A([39]), .B([162]), .Y([163]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10026 (.A([39]), .B([142]), .X([164]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10027 (.A([163]), .B([164]), .Y([165]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10028 (.A([165]), .Y([166]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10029 (.A([167]), .B([143]), .Y([168]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10030 (.A([169]), .B([146]), .Y([170]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10031 (.A([171]), .B([172]), .X([173]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10032 (.A([150]), .B([173]), .Y([174]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10033 (.A([175]), .B([153]), .Y([176]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10034 (.A([170]), .B([176]), .Y([177]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10035 (.A([174]), .B([177]), .X([178]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10036 (.A([178]), .Y([179]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10037 (.A([168]), .B([179]), .Y([180]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10038 (.A([160]), .B([180]), .Y([181]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10039 (.A([181]), .Y([182]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10040 (.A([160]), .B([180]), .X([183]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10041 (.A([181]), .B([183]), .Y([184]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10042 (.A([39]), .B([184]), .Y([185]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10043 (.A([39]), .B([167]), .X([186]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10044 (.A([185]), .B([186]), .Y([187]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10045 (.A([187]), .Y([188]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10046 (.A([189]), .B([143]), .Y([190]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10047 (.A([191]), .B([146]), .Y([192]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10048 (.A([191]), .B([148]), .Y([193]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10049 (.A([194]), .B([153]), .Y([195]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10050 (.A([193]), .B([195]), .Y([196]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10051 (.A([196]), .Y([197]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10052 (.A([192]), .B([197]), .Y([198]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10053 (.A([199]), .B([198]), .X([200]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10054 (.A([200]), .Y([201]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10055 (.A([190]), .B([201]), .Y([202]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10056 (.A([182]), .B([202]), .Y([203]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10057 (.A([203]), .Y([204]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10058 (.A([182]), .B([202]), .X([205]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10059 (.A([203]), .B([205]), .Y([206]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10060 (.A([39]), .B([189]), .X([207]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10061 (.A([39]), .B([206]), .Y([208]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10062 (.A([207]), .B([208]), .Y([209]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10063 (.A([209]), .Y([210]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10064 (.A([211]), .B([143]), .Y([212]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10065 (.A([213]), .B([146]), .Y([214]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10066 (.A([215]), .B([172]), .X([216]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10067 (.A([150]), .B([216]), .Y([217]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10068 (.A([218]), .B([153]), .Y([219]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10069 (.A([214]), .B([219]), .Y([220]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10070 (.A([217]), .B([220]), .X([221]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10071 (.A([221]), .Y([222]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10072 (.A([212]), .B([222]), .Y([223]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10073 (.A([204]), .B([223]), .Y([224]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10074 (.A([224]), .Y([225]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10075 (.A([204]), .B([223]), .X([226]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10076 (.A([224]), .B([226]), .Y([227]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10077 (.A([39]), .B([227]), .Y([228]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10078 (.A([39]), .B([211]), .X([229]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10079 (.A([228]), .B([229]), .Y([230]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10080 (.A([230]), .Y([231]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10081 (.A([232]), .B([143]), .Y([233]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10082 (.A([234]), .B([146]), .Y([235]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10083 (.A([236]), .B([172]), .X([237]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10084 (.A([150]), .B([237]), .Y([238]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10085 (.A([239]), .B([153]), .Y([240]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10086 (.A([235]), .B([240]), .Y([241]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10087 (.A([238]), .B([241]), .X([242]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10088 (.A([242]), .Y([243]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10089 (.A([233]), .B([243]), .Y([244]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10090 (.A([225]), .B([244]), .Y([245]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10091 (.A([245]), .Y([246]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10092 (.A([225]), .B([244]), .X([247]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10093 (.A([245]), .B([247]), .Y([248]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10094 (.A([39]), .B([232]), .X([249]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10095 (.A([39]), .B([248]), .Y([250]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10096 (.A([249]), .B([250]), .Y([251]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10097 (.A([251]), .Y([252]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10098 (.A([253]), .B([254]), .Y([255]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10099 (.A([256]), .B([146]), .Y([257]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10100 (.A([258]), .B([153]), .Y([259]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10101 (.A([258]), .B([148]), .Y([260]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10102 (.A([150]), .B([260]), .Y([261]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10103 (.A([261]), .Y([262]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10104 (.A([263]), .B([264]), .X([265]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10105 (.A([259]), .B([262]), .Y([266]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10106 (.A([257]), .B([265]), .Y([267]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10107 (.A([266]), .B([267]), .X([268]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10108 (.A([268]), .Y([269]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10109 (.A([255]), .B([269]), .Y([270]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10110 (.A([246]), .B([270]), .Y([271]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10111 (.A([271]), .Y([272]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10112 (.A([246]), .B([270]), .X([273]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10113 (.A([271]), .B([273]), .Y([274]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10114 (.A([39]), .B([274]), .Y([275]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10115 (.A([39]), .B([253]), .X([276]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10116 (.A([275]), .B([276]), .Y([277]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10117 (.A([277]), .Y([278]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10118 (.A([279]), .B([254]), .Y([280]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10119 (.A([281]), .B([146]), .Y([282]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10120 (.A([283]), .B([153]), .Y([284]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10121 (.A([283]), .B([148]), .Y([285]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10122 (.A([286]), .B([287]), .Y([288]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10123 (.A([284]), .B([285]), .Y([289]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10124 (.A([199]), .B([289]), .X([290]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10125 (.A([282]), .B([288]), .Y([291]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10126 (.A([290]), .B([291]), .X([292]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10127 (.A([292]), .Y([293]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10128 (.A([280]), .B([293]), .Y([294]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10129 (.A([272]), .B([294]), .Y([295]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10130 (.A([295]), .Y([296]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10131 (.A([272]), .B([294]), .X([297]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10132 (.A([295]), .B([297]), .Y([298]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10133 (.A([39]), .B([298]), .Y([299]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10134 (.A([39]), .B([279]), .X([300]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10135 (.A([299]), .B([300]), .Y([301]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10136 (.A([301]), .Y([302]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10137 (.A([303]), .B([254]), .Y([304]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10138 (.A([305]), .B([146]), .Y([306]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10139 (.A([307]), .B([153]), .Y([308]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10140 (.A([309]), .B([264]), .X([310]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10141 (.A([307]), .B([148]), .Y([311]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10142 (.A([311]), .Y([312]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10143 (.A([150]), .B([308]), .Y([313]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10144 (.A([312]), .B([313]), .X([314]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10145 (.A([306]), .B([310]), .Y([315]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10146 (.A([314]), .B([315]), .X([316]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10147 (.A([316]), .Y([317]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10148 (.A([304]), .B([317]), .Y([318]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10149 (.A([296]), .B([318]), .Y([319]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10150 (.A([319]), .Y([320]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10151 (.A([296]), .B([318]), .X([321]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10152 (.A([319]), .B([321]), .Y([322]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10153 (.A([39]), .B([303]), .X([323]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10154 (.A([39]), .B([322]), .Y([324]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10155 (.A([323]), .B([324]), .Y([325]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10156 (.A([325]), .Y([326]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10157 (.A([327]), .B([254]), .Y([328]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10158 (.A([329]), .B([146]), .Y([330]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10159 (.A([331]), .B([153]), .Y([332]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10160 (.A([145]), .B([287]), .Y([333]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10161 (.A([331]), .B([148]), .Y([334]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10162 (.A([333]), .B([334]), .Y([335]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10163 (.A([199]), .B([335]), .X([336]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10164 (.A([330]), .B([332]), .Y([337]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10165 (.A([336]), .B([337]), .X([338]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10166 (.A([338]), .Y([339]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10167 (.A([328]), .B([339]), .Y([340]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10168 (.A([320]), .B([340]), .Y([341]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10169 (.A([341]), .Y([342]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10170 (.A([320]), .B([340]), .X([343]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10171 (.A([341]), .B([343]), .Y([344]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10172 (.A([39]), .B([344]), .Y([345]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10173 (.A([39]), .B([327]), .X([346]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10174 (.A([345]), .B([346]), .Y([347]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10175 (.A([347]), .Y([348]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10176 (.A([349]), .B([254]), .Y([350]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10177 (.A([350]), .Y([351]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10178 (.A([352]), .B([146]), .Y([353]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10179 (.A([353]), .Y([354]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10180 (.A([355]), .B([153]), .Y([356]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10181 (.A([171]), .B([264]), .X([357]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10182 (.A([355]), .B([148]), .Y([358]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10183 (.A([358]), .Y([359]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10184 (.A([356]), .B([357]), .Y([360]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10185 (.A([359]), .B([360]), .X([361]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10186 (.A([354]), .B([361]), .X([362]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10187 (.A([199]), .B([362]), .X([363]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10188 (.A([351]), .B([363]), .X([364]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10189 (.A([342]), .B([364]), .Y([365]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10190 (.A([365]), .Y([366]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10191 (.A([342]), .B([364]), .X([367]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10192 (.A([365]), .B([367]), .Y([368]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10193 (.A([39]), .B([368]), .Y([369]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10194 (.A([39]), .B([349]), .X([370]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10195 (.A([369]), .B([370]), .Y([371]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10196 (.A([371]), .Y([372]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10197 (.A([373]), .B([254]), .Y([374]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10198 (.A([375]), .B([146]), .Y([376]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10199 (.A([376]), .Y([377]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10200 (.A([378]), .B([153]), .Y([379]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10201 (.A([378]), .B([148]), .Y([380]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10202 (.A([150]), .B([380]), .Y([381]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10203 (.A([191]), .B([287]), .Y([382]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10204 (.A([379]), .B([382]), .Y([383]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10205 (.A([381]), .B([383]), .X([384]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10206 (.A([384]), .Y([385]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10207 (.A([374]), .B([385]), .Y([386]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10208 (.A([377]), .B([386]), .X([387]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10209 (.A([366]), .B([387]), .Y([388]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10210 (.A([388]), .Y([389]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10211 (.A([366]), .B([387]), .X([390]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10212 (.A([388]), .B([390]), .Y([391]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10213 (.A([39]), .B([391]), .Y([392]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10214 (.A([39]), .B([373]), .X([393]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10215 (.A([392]), .B([393]), .Y([394]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10216 (.A([394]), .Y([395]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10217 (.A([396]), .B([254]), .Y([397]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10218 (.A([398]), .B([146]), .Y([399]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10219 (.A([400]), .B([148]), .Y([401]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10220 (.A([215]), .B([264]), .X([402]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10221 (.A([401]), .B([402]), .Y([403]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10222 (.A([199]), .B([403]), .X([404]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10223 (.A([400]), .B([153]), .Y([405]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10224 (.A([399]), .B([405]), .Y([406]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10225 (.A([404]), .B([406]), .X([407]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10226 (.A([407]), .Y([408]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10227 (.A([397]), .B([408]), .Y([409]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10228 (.A([389]), .B([409]), .Y([410]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10229 (.A([389]), .B([409]), .X([411]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10230 (.A([410]), .B([411]), .Y([412]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10231 (.A([39]), .B([412]), .Y([413]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10232 (.A([39]), .B([396]), .X([414]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10233 (.A([413]), .B([414]), .Y([415]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10234 (.A([415]), .Y([416]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10235 (.A([417]), .B([254]), .Y([418]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10236 (.A([419]), .B([146]), .Y([420]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10237 (.A([421]), .B([153]), .Y([422]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10238 (.A([236]), .B([264]), .X([423]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10239 (.A([421]), .B([148]), .Y([424]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10240 (.A([420]), .B([423]), .Y([425]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10241 (.A([422]), .B([424]), .Y([426]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10242 (.A([199]), .B([426]), .X([427]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10243 (.A([425]), .B([427]), .X([428]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10244 (.A([428]), .Y([429]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10245 (.A([418]), .B([429]), .Y([430]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10246 (.A([410]), .B([430]), .X([431]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10247 (.A([410]), .B([430]), .Y([432]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10248 (.A([433]), .B([417]), .Y([434]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10249 (.A([431]), .B([432]), .Y([435]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10250 (.A([39]), .B([435]), .Y([436]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10251 (.A([434]), .B([436]), .Y([437]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10252 (.A([433]), .B([438]), .Y([439]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10253 (.A([39]), .B([440]), .Y([441]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10254 (.A([439]), .B([441]), .Y([442]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10255 (.A([433]), .B([443]), .Y([444]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10256 (.A([39]), .B([445]), .Y([446]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10257 (.A([444]), .B([446]), .Y([447]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10258 (.A([433]), .B([448]), .Y([449]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10259 (.A([39]), .B([450]), .Y([451]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10260 (.A([449]), .B([451]), .Y([452]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10261 (.A([453]), .B([454]), .X([455]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10262 (.A([453]), .B([456]), .Y([457]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10263 (.A([60]), .B([454]), .Y([458]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10264 (.A([459]), .B([458]), .Y([460]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10265 (.A([457]), .B([460]), .Y([461]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10266 (.A([462]), .B([461]), .X([463]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10267 (.A([462]), .B([145]), .Y([464]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10268 (.A([463]), .B([464]), .Y([465]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10269 (.A([466]), .B([465]), .Y([467]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10270 (.A([468]), .B([469]), .X([470]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10271 (.A([470]), .Y([471]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10272 (.A([472]), .B([455]), .Y([473]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10273 (.A([474]), .B([469]), .Y([475]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10274 (.A([476]), .B([473]), .Y([477]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10275 (.A([475]), .B([477]), .X([478]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10276 (.A([467]), .B([478]), .Y([479]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10277 (.A([471]), .B([479]), .X([480]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10278 (.A([481]), .B([482]), .Y([483]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10279 (.A([484]), .B([483]), .Y([485]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10280 (.A([472]), .B([485]), .Y([486]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10281 (.A([476]), .B([486]), .Y([487]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10282 (.A([488]), .B([489]), .X([490]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10283 (.A([490]), .Y([491]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10284 (.A([469]), .B([490]), .Y([492]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10285 (.A([492]), .Y([493]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10286 (.A([494]), .B([493]), .Y([495]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10287 (.A([496]), .B([495]), .X([497]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10288 (.A([487]), .B([497]), .X([498]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10289 (.A([236]), .B([490]), .X([499]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10290 (.A([419]), .B([490]), .Y([500]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10291 (.A([501]), .B([500]), .X([502]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10292 (.A([499]), .B([502]), .Y([503]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10293 (.A([234]), .B([487]), .Y([504]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10294 (.A([492]), .B([504]), .X([505]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10295 (.A([498]), .B([505]), .Y([506]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10296 (.A([503]), .B([506]), .X([507]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10297 (.A([508]), .B([469]), .X([509]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10298 (.A([462]), .B([286]), .Y([510]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10299 (.A([511]), .B([485]), .X([512]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10300 (.A([145]), .B([169]), .X([513]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10301 (.A([191]), .B([213]), .X([514]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10302 (.A([513]), .B([514]), .X([515]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10303 (.A([234]), .B([516]), .X([517]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10304 (.A([286]), .B([518]), .X([519]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10305 (.A([517]), .B([519]), .X([520]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10306 (.A([515]), .B([520]), .X([521]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10307 (.A([462]), .B([521]), .X([522]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10308 (.A([522]), .Y([523]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10309 (.A([512]), .B([523]), .Y([524]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10310 (.A([510]), .B([524]), .Y([525]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10311 (.A([466]), .B([525]), .Y([526]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10312 (.A([509]), .B([526]), .Y([527]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10313 (.A([490]), .B([527]), .Y([528]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10314 (.A([490]), .B([521]), .X([529]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10315 (.A([472]), .B([512]), .Y([530]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10316 (.A([531]), .B([476]), .Y([532]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10317 (.A([492]), .B([532]), .X([533]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10318 (.A([533]), .Y([534]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10319 (.A([530]), .B([534]), .Y([535]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10320 (.A([529]), .B([535]), .Y([536]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10321 (.A([536]), .Y([537]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10322 (.A([528]), .B([537]), .Y([538]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10323 (.A([539]), .B([491]), .Y([540]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10324 (.A([540]), .Y([541]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10325 (.A([542]), .B([540]), .Y([543]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10326 (.A([544]), .B([539]), .X([545]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10327 (.A([546]), .B([545]), .X([547]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10328 (.A([547]), .Y([548]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10329 (.A([543]), .B([547]), .Y([549]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10330 (.A([550]), .B([549]), .X([551]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10331 (.A([60]), .B([552]), .Y([553]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10332 (.A([554]), .B([44]), .Y([555]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10333 (.A([554]), .B([553]), .X([556]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10334 (.A([555]), .B([556]), .Y([557]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10335 (.A([462]), .B([557]), .X([558]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10336 (.A([462]), .B([263]), .Y([559]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10337 (.A([558]), .B([559]), .Y([560]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10338 (.A([548]), .B([560]), .Y([561]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10339 (.A([562]), .B([472]), .Y([563]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10340 (.A([563]), .Y([564]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10341 (.A([561]), .B([564]), .Y([565]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10342 (.A([542]), .B([565]), .X([566]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10343 (.A([567]), .B([469]), .X([568]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10344 (.A([540]), .B([568]), .Y([569]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10345 (.A([569]), .Y([570]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10346 (.A([566]), .B([570]), .Y([571]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10347 (.A([551]), .B([571]), .Y([572]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10348 (.A([462]), .B([554]), .X([573]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10349 (.A([552]), .B([573]), .X([574]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10350 (.A([547]), .B([574]), .X([575]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10351 (.A([564]), .B([575]), .Y([576]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10352 (.A([577]), .B([469]), .Y([578]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10353 (.A([578]), .Y([579]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10354 (.A([576]), .B([579]), .Y([580]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10355 (.A([541]), .B([580]), .X([581]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10356 (.A([572]), .B([581]), .Y([582]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10357 (.A([433]), .B([583]), .Y([584]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10358 (.A([585]), .B([584]), .Y([586]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10359 (.A([587]), .B([588]), .X([589]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10360 (.A([590]), .B([588]), .Y([591]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10361 (.A([589]), .B([591]), .Y([592]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10362 (.A([593]), .B([592]), .Y([594]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10363 (.A([595]), .B([588]), .X([596]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10364 (.A([597]), .B([588]), .Y([598]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10365 (.A([596]), .B([598]), .Y([599]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10366 (.A([600]), .B([599]), .Y([601]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10367 (.A([594]), .B([601]), .Y([602]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10368 (.A([603]), .B([602]), .Y([604]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10369 (.A([605]), .B([606]), .X([607]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10370 (.A([608]), .B([609]), .X([610]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10371 (.A([611]), .B([610]), .X([612]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10372 (.A([607]), .B([612]), .Y([613]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10373 (.A([614]), .B([615]), .X([616]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10374 (.A([617]), .B([616]), .Y([618]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10375 (.A([613]), .B([618]), .X([619]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10376 (.A([469]), .B([150]), .Y([620]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10377 (.A([488]), .B([621]), .X([622]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10378 (.A([614]), .B([623]), .X([624]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10379 (.A([622]), .B([624]), .Y([625]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10380 (.A([620]), .B([625]), .X([626]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10381 (.A([488]), .B([623]), .X([627]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10382 (.A([627]), .Y([628]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10383 (.A([629]), .B([627]), .Y([630]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10384 (.A([605]), .B([631]), .X([632]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10385 (.A([632]), .Y([633]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10386 (.A([634]), .B([630]), .X([635]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10387 (.A([626]), .B([633]), .X([636]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10388 (.A([635]), .B([636]), .X([637]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10389 (.A([637]), .Y([638]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10390 (.A([605]), .B([639]), .X([640]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10391 (.A([641]), .B([642]), .X([643]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10392 (.A([614]), .B([643]), .X([644]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10393 (.A([640]), .B([644]), .Y([645]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10394 (.A([614]), .B([610]), .X([646]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10395 (.A([605]), .B([610]), .X([647]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10396 (.A([646]), .B([647]), .Y([648]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10397 (.A([645]), .B([648]), .X([649]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10398 (.A([650]), .B([649]), .X([651]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10399 (.A([619]), .B([651]), .X([652]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10400 (.A([637]), .B([652]), .X([653]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10401 (.A([614]), .B([654]), .X([655]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10402 (.A([655]), .Y([656]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10403 (.A([605]), .B([643]), .X([657]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10404 (.A([264]), .B([657]), .Y([658]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10405 (.A([656]), .B([658]), .X([659]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10406 (.A([488]), .B([643]), .X([660]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10407 (.A([660]), .Y([661]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10408 (.A([488]), .B([639]), .X([662]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10409 (.A([660]), .B([662]), .Y([663]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10410 (.A([491]), .B([663]), .X([664]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10411 (.A([659]), .B([664]), .X([665]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10412 (.A([666]), .B([614]), .X([667]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10413 (.A([488]), .B([606]), .X([668]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10414 (.A([667]), .B([668]), .Y([669]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10415 (.A([148]), .B([669]), .X([670]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10416 (.A([603]), .B([670]), .X([671]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10417 (.A([665]), .B([671]), .X([672]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10418 (.A([653]), .B([672]), .X([673]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10419 (.A([673]), .Y([674]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10420 (.A([675]), .B([674]), .Y([676]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10421 (.A([516]), .B([653]), .Y([677]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10422 (.A([678]), .B([665]), .Y([679]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10423 (.A([256]), .B([669]), .Y([680]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10424 (.A([681]), .B([680]), .Y([682]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10425 (.A([682]), .Y([683]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10426 (.A([679]), .B([683]), .Y([684]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10427 (.A([684]), .Y([685]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10428 (.A([677]), .B([685]), .Y([686]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10429 (.A([686]), .Y([687]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10430 (.A([676]), .B([687]), .Y([688]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10431 (.A([688]), .Y([689]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10432 (.A([604]), .B([689]), .Y([84]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10433 (.A([690]), .B([691]), .Y([692]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10434 (.A([488]), .B([610]), .X([693]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10435 (.A([694]), .B([693]), .Y([695]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10436 (.A([695]), .Y([696]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10437 (.A([697]), .B([695]), .X([698]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10438 (.A([39]), .B([692]), .Y([699]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10439 (.A([698]), .B([699]), .X([700]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10440 (.A([700]), .Y([701]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10441 (.A([84]), .B([701]), .Y([702]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10442 (.A([678]), .B([700]), .Y([703]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10443 (.A([702]), .B([703]), .Y([704]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10444 (.A([705]), .B([588]), .Y([706]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10445 (.A([707]), .B([588]), .X([708]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10446 (.A([706]), .B([708]), .Y([709]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10447 (.A([600]), .B([709]), .Y([710]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10448 (.A([711]), .B([482]), .X([712]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10449 (.A([712]), .Y([713]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10450 (.A([714]), .B([715]), .X([716]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10451 (.A([710]), .B([716]), .Y([717]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10452 (.A([713]), .B([717]), .X([718]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10453 (.A([719]), .B([718]), .X([720]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10454 (.A([721]), .B([674]), .Y([722]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10455 (.A([286]), .B([653]), .Y([723]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10456 (.A([724]), .B([665]), .Y([725]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10457 (.A([281]), .B([669]), .Y([726]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10458 (.A([725]), .B([726]), .Y([727]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10459 (.A([722]), .B([723]), .Y([728]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10460 (.A([729]), .B([728]), .X([730]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10461 (.A([727]), .B([730]), .X([731]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10462 (.A([731]), .Y([732]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10463 (.A([720]), .B([732]), .Y([85]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10464 (.A([701]), .B([85]), .Y([733]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10465 (.A([724]), .B([700]), .Y([734]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10466 (.A([733]), .B([734]), .Y([735]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10467 (.A([736]), .B([737]), .Y([738]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10468 (.A([739]), .B([588]), .Y([740]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10469 (.A([738]), .B([740]), .Y([741]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10470 (.A([593]), .B([741]), .X([742]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10471 (.A([743]), .B([482]), .X([744]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10472 (.A([744]), .Y([745]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10473 (.A([746]), .B([715]), .X([747]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10474 (.A([742]), .B([747]), .Y([748]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10475 (.A([745]), .B([748]), .X([749]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10476 (.A([719]), .B([749]), .X([750]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10477 (.A([138]), .B([674]), .Y([751]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10478 (.A([518]), .B([653]), .Y([752]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10479 (.A([753]), .B([665]), .Y([754]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10480 (.A([305]), .B([669]), .Y([755]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10481 (.A([754]), .B([755]), .Y([756]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10482 (.A([124]), .B([756]), .X([757]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10483 (.A([757]), .Y([758]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10484 (.A([752]), .B([758]), .Y([759]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10485 (.A([759]), .Y([760]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10486 (.A([751]), .B([760]), .Y([761]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10487 (.A([761]), .Y([762]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10488 (.A([750]), .B([762]), .Y([86]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10489 (.A([701]), .B([86]), .Y([763]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10490 (.A([753]), .B([700]), .Y([764]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10491 (.A([763]), .B([764]), .Y([765]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10492 (.A([766]), .B([737]), .Y([767]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10493 (.A([768]), .B([588]), .Y([769]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10494 (.A([767]), .B([769]), .Y([770]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10495 (.A([593]), .B([770]), .X([771]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10496 (.A([772]), .B([715]), .X([773]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10497 (.A([773]), .Y([774]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10498 (.A([775]), .B([482]), .X([776]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10499 (.A([771]), .B([776]), .Y([777]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10500 (.A([774]), .B([777]), .X([778]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10501 (.A([719]), .B([778]), .X([779]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10502 (.A([142]), .B([674]), .Y([780]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10503 (.A([145]), .B([653]), .Y([781]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10504 (.A([152]), .B([665]), .Y([782]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10505 (.A([329]), .B([669]), .Y([783]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10506 (.A([149]), .B([783]), .Y([784]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10507 (.A([784]), .Y([785]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10508 (.A([782]), .B([785]), .Y([786]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10509 (.A([786]), .Y([787]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10510 (.A([781]), .B([787]), .Y([788]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10511 (.A([788]), .Y([789]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10512 (.A([780]), .B([789]), .Y([790]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10513 (.A([790]), .Y([791]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10514 (.A([779]), .B([791]), .Y([87]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10515 (.A([152]), .B([700]), .Y([792]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10516 (.A([701]), .B([87]), .Y([793]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10517 (.A([792]), .B([793]), .Y([794]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10518 (.A([795]), .B([737]), .Y([796]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10519 (.A([797]), .B([588]), .Y([798]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10520 (.A([796]), .B([798]), .Y([799]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10521 (.A([593]), .B([799]), .X([800]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10522 (.A([801]), .B([482]), .X([802]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10523 (.A([802]), .Y([803]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10524 (.A([804]), .B([715]), .X([805]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10525 (.A([800]), .B([805]), .Y([806]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10526 (.A([803]), .B([806]), .X([807]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10527 (.A([719]), .B([807]), .X([808]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10528 (.A([167]), .B([674]), .Y([809]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10529 (.A([169]), .B([653]), .Y([810]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10530 (.A([175]), .B([665]), .Y([811]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10531 (.A([352]), .B([669]), .Y([812]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10532 (.A([173]), .B([812]), .Y([813]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10533 (.A([813]), .Y([814]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10534 (.A([811]), .B([814]), .Y([815]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10535 (.A([815]), .Y([816]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10536 (.A([810]), .B([816]), .Y([817]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10537 (.A([817]), .Y([818]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10538 (.A([809]), .B([818]), .Y([819]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10539 (.A([819]), .Y([820]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10540 (.A([808]), .B([820]), .Y([88]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10541 (.A([701]), .B([88]), .Y([821]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10542 (.A([175]), .B([700]), .Y([822]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10543 (.A([821]), .B([822]), .Y([823]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10544 (.A([824]), .B([737]), .Y([825]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10545 (.A([826]), .B([588]), .Y([827]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10546 (.A([825]), .B([827]), .Y([828]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10547 (.A([593]), .B([828]), .X([829]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10548 (.A([830]), .B([482]), .X([831]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10549 (.A([831]), .Y([832]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10550 (.A([833]), .B([715]), .X([834]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10551 (.A([829]), .B([834]), .Y([835]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10552 (.A([832]), .B([835]), .X([836]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10553 (.A([719]), .B([836]), .X([837]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10554 (.A([189]), .B([674]), .Y([838]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10555 (.A([191]), .B([653]), .Y([839]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10556 (.A([194]), .B([665]), .Y([840]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10557 (.A([375]), .B([669]), .Y([841]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10558 (.A([193]), .B([841]), .Y([842]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10559 (.A([842]), .Y([843]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10560 (.A([840]), .B([843]), .Y([844]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10561 (.A([844]), .Y([845]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10562 (.A([839]), .B([845]), .Y([846]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10563 (.A([846]), .Y([847]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10564 (.A([838]), .B([847]), .Y([848]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10565 (.A([848]), .Y([849]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10566 (.A([837]), .B([849]), .Y([89]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10567 (.A([701]), .B([89]), .Y([850]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10568 (.A([194]), .B([700]), .Y([851]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10569 (.A([850]), .B([851]), .Y([852]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10570 (.A([853]), .B([737]), .Y([854]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10571 (.A([855]), .B([588]), .Y([856]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10572 (.A([854]), .B([856]), .Y([857]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10573 (.A([593]), .B([857]), .X([858]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10574 (.A([859]), .B([482]), .X([860]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10575 (.A([860]), .Y([861]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10576 (.A([862]), .B([715]), .X([863]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10577 (.A([858]), .B([863]), .Y([864]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10578 (.A([861]), .B([864]), .X([865]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10579 (.A([719]), .B([865]), .X([866]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10580 (.A([211]), .B([674]), .Y([867]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10581 (.A([213]), .B([653]), .Y([868]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10582 (.A([218]), .B([665]), .Y([869]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10583 (.A([398]), .B([669]), .Y([870]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10584 (.A([216]), .B([870]), .Y([871]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10585 (.A([871]), .Y([872]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10586 (.A([869]), .B([872]), .Y([873]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10587 (.A([873]), .Y([874]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10588 (.A([868]), .B([874]), .Y([875]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10589 (.A([875]), .Y([876]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10590 (.A([867]), .B([876]), .Y([877]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10591 (.A([877]), .Y([878]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10592 (.A([866]), .B([878]), .Y([90]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10593 (.A([218]), .B([700]), .Y([879]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10594 (.A([701]), .B([90]), .Y([880]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10595 (.A([879]), .B([880]), .Y([881]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10596 (.A([882]), .B([737]), .Y([883]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10597 (.A([884]), .B([588]), .Y([885]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10598 (.A([883]), .B([885]), .Y([886]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10599 (.A([593]), .B([886]), .X([887]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10600 (.A([888]), .B([715]), .X([889]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10601 (.A([889]), .Y([890]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10602 (.A([891]), .B([482]), .X([892]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10603 (.A([887]), .B([892]), .Y([893]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10604 (.A([890]), .B([893]), .X([894]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10605 (.A([719]), .B([894]), .X([895]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10606 (.A([232]), .B([674]), .Y([896]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10607 (.A([234]), .B([653]), .Y([897]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10608 (.A([239]), .B([665]), .Y([898]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10609 (.A([419]), .B([669]), .Y([899]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10610 (.A([899]), .Y([900]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10611 (.A([237]), .B([895]), .Y([901]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10612 (.A([897]), .B([898]), .Y([902]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10613 (.A([902]), .Y([903]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10614 (.A([896]), .B([903]), .Y([904]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10615 (.A([900]), .B([904]), .X([905]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10616 (.A([901]), .B([905]), .X([91]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10617 (.A([701]), .B([91]), .Y([906]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10618 (.A([239]), .B([700]), .Y([907]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10619 (.A([906]), .B([907]), .Y([908]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10620 (.A([253]), .B([674]), .Y([909]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10621 (.A([256]), .B([651]), .Y([910]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10622 (.A([638]), .B([910]), .Y([911]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10623 (.A([719]), .B([260]), .Y([912]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10624 (.A([258]), .B([664]), .Y([913]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10625 (.A([516]), .B([659]), .Y([914]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10626 (.A([913]), .B([914]), .Y([915]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10627 (.A([912]), .B([915]), .X([916]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10628 (.A([911]), .B([916]), .X([917]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10629 (.A([917]), .Y([918]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10630 (.A([909]), .B([918]), .Y([92]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10631 (.A([258]), .B([700]), .Y([919]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10632 (.A([701]), .B([92]), .Y([920]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10633 (.A([919]), .B([920]), .Y([921]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10634 (.A([279]), .B([674]), .Y([922]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10635 (.A([281]), .B([651]), .Y([923]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10636 (.A([283]), .B([664]), .Y([924]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10637 (.A([286]), .B([659]), .Y([925]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10638 (.A([285]), .B([925]), .Y([926]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10639 (.A([923]), .B([924]), .Y([927]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10640 (.A([926]), .B([927]), .X([928]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10641 (.A([928]), .Y([929]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10642 (.A([922]), .B([929]), .Y([93]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10643 (.A([283]), .B([700]), .Y([930]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10644 (.A([701]), .B([93]), .Y([931]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10645 (.A([930]), .B([931]), .Y([932]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10646 (.A([303]), .B([674]), .Y([933]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10647 (.A([305]), .B([651]), .Y([934]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10648 (.A([518]), .B([659]), .Y([935]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10649 (.A([307]), .B([664]), .Y([936]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10650 (.A([934]), .B([936]), .Y([937]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10651 (.A([311]), .B([935]), .Y([938]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10652 (.A([937]), .B([938]), .X([939]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10653 (.A([939]), .Y([940]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10654 (.A([933]), .B([940]), .Y([94]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10655 (.A([307]), .B([700]), .Y([941]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10656 (.A([701]), .B([94]), .Y([942]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10657 (.A([941]), .B([942]), .Y([943]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10658 (.A([327]), .B([674]), .Y([944]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10659 (.A([329]), .B([651]), .Y([945]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10660 (.A([145]), .B([659]), .Y([946]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10661 (.A([331]), .B([664]), .Y([947]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10662 (.A([334]), .B([947]), .Y([948]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10663 (.A([945]), .B([946]), .Y([949]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10664 (.A([948]), .B([949]), .X([950]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10665 (.A([950]), .Y([951]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10666 (.A([944]), .B([951]), .Y([95]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10667 (.A([701]), .B([95]), .Y([952]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10668 (.A([331]), .B([700]), .Y([953]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10669 (.A([952]), .B([953]), .Y([954]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10670 (.A([349]), .B([674]), .Y([955]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10671 (.A([352]), .B([651]), .Y([956]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10672 (.A([169]), .B([659]), .Y([957]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10673 (.A([355]), .B([664]), .Y([958]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10674 (.A([956]), .B([958]), .Y([959]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10675 (.A([358]), .B([957]), .Y([960]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10676 (.A([959]), .B([960]), .X([961]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10677 (.A([961]), .Y([962]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10678 (.A([955]), .B([962]), .Y([96]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10679 (.A([701]), .B([96]), .Y([963]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10680 (.A([355]), .B([700]), .Y([964]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10681 (.A([963]), .B([964]), .Y([965]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10682 (.A([373]), .B([674]), .Y([966]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10683 (.A([375]), .B([651]), .Y([967]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10684 (.A([378]), .B([664]), .Y([968]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10685 (.A([191]), .B([659]), .Y([969]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10686 (.A([380]), .B([969]), .Y([970]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10687 (.A([967]), .B([968]), .Y([971]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10688 (.A([970]), .B([971]), .X([972]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10689 (.A([972]), .Y([973]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10690 (.A([966]), .B([973]), .Y([97]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10691 (.A([701]), .B([97]), .Y([974]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10692 (.A([378]), .B([700]), .Y([975]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10693 (.A([974]), .B([975]), .Y([976]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10694 (.A([396]), .B([674]), .Y([977]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10695 (.A([398]), .B([651]), .Y([978]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10696 (.A([978]), .Y([979]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10697 (.A([213]), .B([659]), .Y([980]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10698 (.A([980]), .Y([981]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10699 (.A([400]), .B([664]), .Y([982]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10700 (.A([401]), .B([982]), .Y([983]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10701 (.A([981]), .B([983]), .X([984]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10702 (.A([979]), .B([984]), .X([985]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10703 (.A([985]), .Y([986]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10704 (.A([977]), .B([986]), .Y([98]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10705 (.A([701]), .B([98]), .Y([987]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10706 (.A([400]), .B([700]), .Y([988]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10707 (.A([987]), .B([988]), .Y([989]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10708 (.A([417]), .B([674]), .Y([990]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10709 (.A([419]), .B([651]), .Y([991]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10710 (.A([234]), .B([659]), .Y([992]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10711 (.A([421]), .B([664]), .Y([993]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10712 (.A([424]), .B([993]), .Y([994]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10713 (.A([991]), .B([992]), .Y([995]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10714 (.A([994]), .B([995]), .X([996]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10715 (.A([996]), .Y([997]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10716 (.A([990]), .B([997]), .Y([99]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10717 (.A([701]), .B([99]), .Y([998]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10718 (.A([421]), .B([700]), .Y([999]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10719 (.A([998]), .B([999]), .Y([1000]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10720 (.A([39]), .B([695]), .Y([1001]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10721 (.A([1002]), .B([1001]), .X([1003]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10722 (.A([1003]), .Y([1004]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10723 (.A([567]), .B([1003]), .X([1005]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10724 (.A([1006]), .B([1003]), .Y([1007]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10725 (.A([1005]), .B([1007]), .Y([1008]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10726 (.A([508]), .B([1003]), .X([1009]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10727 (.A([1010]), .B([1003]), .Y([1011]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10728 (.A([1009]), .B([1011]), .Y([1012]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10729 (.A([1013]), .B([1003]), .Y([1014]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10730 (.A([1015]), .B([1003]), .X([1016]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10731 (.A([1014]), .B([1016]), .Y([1017]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10732 (.A([468]), .B([1003]), .X([1018]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10733 (.A([1019]), .B([1003]), .Y([1020]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10734 (.A([1018]), .B([1020]), .Y([1021]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10735 (.A([352]), .B([1004]), .Y([1022]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10736 (.A([1023]), .B([1003]), .Y([1024]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10737 (.A([1022]), .B([1024]), .Y([1025]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10738 (.A([1026]), .B([1003]), .Y([1027]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10739 (.A([1028]), .B([1003]), .X([1029]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10740 (.A([1027]), .B([1029]), .Y([1030]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10741 (.A([1031]), .B([1003]), .Y([1032]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10742 (.A([1033]), .B([1003]), .X([1034]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10743 (.A([1032]), .B([1034]), .Y([1035]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10744 (.A([1036]), .B([1003]), .Y([1037]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10745 (.A([419]), .B([1004]), .Y([1038]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10746 (.A([1037]), .B([1038]), .Y([1039]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10747 (.A([1040]), .B([1041]), .Y([1042]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10748 (.A([1043]), .B([1042]), .Y([1044]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10749 (.A([1044]), .Y([1045]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10750 (.A([1046]), .B([1047]), .X([1048]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10751 (.A([1049]), .B([1050]), .X([1051]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10752 (.A([1052]), .B([1051]), .X([1053]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10753 (.A([1048]), .B([1053]), .Y([1054]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10754 (.A([1055]), .B([1056]), .X([1057]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10755 (.A([1058]), .B([1057]), .X([1059]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10756 (.A([1059]), .Y([1060]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10757 (.A([1061]), .B([1062]), .X([1063]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10758 (.A([1064]), .B([1063]), .Y([1065]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10759 (.A([1066]), .B([1065]), .X([1067]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10760 (.A([1060]), .B([1067]), .X([1068]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10761 (.A([1069]), .B([1062]), .Y([1070]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10762 (.A([1070]), .Y([1071]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10763 (.A([1072]), .B([1073]), .Y([1074]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10764 (.A([1071]), .B([1074]), .Y([1075]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10765 (.A([1047]), .B([1076]), .X([1077]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10766 (.A([1077]), .Y([1078]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10767 (.A([1075]), .B([1077]), .Y([1079]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10768 (.A([1068]), .B([1079]), .X([1080]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10769 (.A([1054]), .B([1080]), .X([1081]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10770 (.A([1045]), .B([1081]), .X([1082]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10771 (.A([1083]), .B([1047]), .X([1084]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10772 (.A([1085]), .B([1084]), .Y([1086]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10773 (.A([1087]), .B([1088]), .X([1089]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10774 (.A([1057]), .B([1089]), .X([1090]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10775 (.A([1052]), .B([1089]), .X([1091]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10776 (.A([1090]), .B([1091]), .Y([1092]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10777 (.A([1086]), .B([1092]), .X([1093]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10778 (.A([1094]), .B([1095]), .X([1096]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10779 (.A([1097]), .B([1041]), .X([1098]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10780 (.A([1056]), .B([1098]), .X([1099]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10781 (.A([1096]), .B([1099]), .Y([1100]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10782 (.A([1101]), .B([1057]), .X([1102]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10783 (.A([1095]), .B([1070]), .Y([1103]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10784 (.A([1094]), .B([1103]), .Y([1104]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10785 (.A([1046]), .B([1057]), .X([1105]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10786 (.A([1104]), .B([1105]), .Y([1106]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10787 (.A([1106]), .Y([1107]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10788 (.A([1102]), .B([1107]), .Y([1108]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10789 (.A([1100]), .B([1108]), .X([1109]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10790 (.A([1093]), .B([1109]), .X([1110]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10791 (.A([1082]), .B([1110]), .X([1111]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10792 (.A([264]), .B([692]), .Y([1112]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10793 (.A([1113]), .B([660]), .Y([1114]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10794 (.A([1115]), .B([1114]), .X([1116]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10795 (.A([1112]), .B([1116]), .X([1117]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10796 (.A([646]), .B([655]), .Y([1118]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10797 (.A([1119]), .B([1118]), .X([1120]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10798 (.A([491]), .B([1120]), .X([1121]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10799 (.A([1121]), .Y([1122]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10800 (.A([1123]), .B([691]), .Y([1124]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10801 (.A([1125]), .B([1126]), .Y([1127]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10802 (.A([1127]), .Y([1128]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10803 (.A([1124]), .B([1128]), .Y([1129]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10804 (.A([617]), .B([1130]), .Y([1131]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10805 (.A([1132]), .B([1133]), .Y([1134]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10806 (.A([1131]), .B([1134]), .X([1135]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10807 (.A([1129]), .B([1135]), .X([1136]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10808 (.A([1121]), .B([1136]), .X([1137]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10809 (.A([1117]), .B([1137]), .X([1138]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10810 (.A([469]), .B([622]), .Y([1139]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10811 (.A([630]), .B([1139]), .X([1140]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10812 (.A([1141]), .B([1140]), .X([1142]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10813 (.A([1143]), .B([1144]), .X([1145]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10814 (.A([1142]), .B([1145]), .X([1146]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10815 (.A([645]), .B([695]), .X([1147]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10816 (.A([647]), .B([657]), .Y([1148]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10817 (.A([624]), .B([632]), .Y([1149]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10818 (.A([1148]), .B([1149]), .X([1150]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10819 (.A([1147]), .B([1150]), .X([1151]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10820 (.A([662]), .B([668]), .Y([1152]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10821 (.A([614]), .B([1153]), .X([1154]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10822 (.A([1154]), .Y([1155]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10823 (.A([614]), .B([621]), .X([1156]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10824 (.A([1156]), .Y([1157]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10825 (.A([1154]), .B([1156]), .Y([1158]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10826 (.A([1152]), .B([1158]), .X([1159]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10827 (.A([1160]), .B([1161]), .Y([1162]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10828 (.A([613]), .B([1162]), .X([1163]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10829 (.A([1159]), .B([1163]), .X([1164]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10830 (.A([1151]), .B([1164]), .X([1165]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10831 (.A([1146]), .B([1165]), .X([1166]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10832 (.A([1138]), .B([1166]), .X([1167]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10833 (.A([39]), .B([1167]), .Y([1168]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10834 (.A([1168]), .Y([1169]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10835 (.A([1051]), .B([1057]), .X([1170]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10836 (.A([1040]), .B([1057]), .X([1171]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10837 (.A([1111]), .B([1169]), .Y([1172]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10838 (.A([1172]), .Y([1173]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10839 (.A([1174]), .B([1063]), .X([1175]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10840 (.A([1175]), .Y([1176]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10841 (.A([1100]), .B([1176]), .X([1177]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10842 (.A([1060]), .B([1177]), .X([1178]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10843 (.A([1077]), .B([1090]), .Y([1179]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10844 (.A([1178]), .B([1179]), .X([1180]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10845 (.A([472]), .B([1180]), .Y([1181]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10846 (.A([612]), .B([668]), .Y([1182]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10847 (.A([1148]), .B([1182]), .X([1183]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10848 (.A([172]), .B([1184]), .X([1185]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10849 (.A([1156]), .B([1185]), .Y([1186]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10850 (.A([1160]), .B([150]), .Y([1187]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10851 (.A([1161]), .B([1188]), .Y([1189]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10852 (.A([1187]), .B([1189]), .X([1190]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10853 (.A([1186]), .B([1190]), .X([1191]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10854 (.A([1183]), .B([1191]), .X([1192]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10855 (.A([1193]), .B([550]), .X([1194]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10856 (.A([1194]), .Y([1195]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10857 (.A([1196]), .B([1194]), .X([1197]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10858 (.A([640]), .B([1197]), .X([1198]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10859 (.A([1124]), .B([1198]), .Y([1199]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10860 (.A([1200]), .B([1201]), .Y([1202]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10861 (.A([1199]), .B([1202]), .X([1203]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10862 (.A([1130]), .B([622]), .Y([1204]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10863 (.A([1155]), .B([1204]), .X([1205]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10864 (.A([629]), .B([694]), .Y([1206]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10865 (.A([1133]), .B([644]), .Y([1207]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10866 (.A([1206]), .B([1207]), .X([1208]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10867 (.A([1205]), .B([1208]), .X([1209]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10868 (.A([1203]), .B([1209]), .X([1210]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10869 (.A([1121]), .B([1210]), .X([1211]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10870 (.A([1192]), .B([1211]), .X([1212]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10871 (.A([1212]), .Y([1213]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10872 (.A([1181]), .B([1213]), .Y([1214]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10873 (.A([1173]), .B([1214]), .Y([1215]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10874 (.A([1216]), .B([1172]), .Y([1217]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10875 (.A([1215]), .B([1217]), .Y([1218]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10876 (.A([1219]), .B([1091]), .Y([1220]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10877 (.A([1094]), .B([1064]), .X([1221]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10878 (.A([1048]), .B([1221]), .Y([1222]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10879 (.A([1222]), .Y([1223]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10880 (.A([1106]), .B([1176]), .X([1224]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10881 (.A([1222]), .B([1224]), .X([1225]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10882 (.A([1220]), .B([1225]), .X([1226]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10883 (.A([472]), .B([1226]), .Y([1227]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10884 (.A([438]), .B([443]), .X([1228]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10885 (.A([1228]), .Y([1229]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10886 (.A([1230]), .B([1229]), .Y([1231]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10887 (.A([438]), .B([1232]), .X([1233]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10888 (.A([1233]), .Y([1234]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10889 (.A([1235]), .B([1234]), .Y([1236]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10890 (.A([1231]), .B([1236]), .Y([1237]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10891 (.A([1238]), .B([1232]), .X([1239]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10892 (.A([1240]), .B([1239]), .X([1241]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10893 (.A([443]), .B([1238]), .X([1242]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10894 (.A([1243]), .B([1242]), .X([1244]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10895 (.A([1241]), .B([1244]), .Y([1245]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10896 (.A([1237]), .B([1245]), .X([1246]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10897 (.A([1247]), .B([1246]), .Y([1248]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10898 (.A([1249]), .B([1229]), .Y([1250]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10899 (.A([1251]), .B([1234]), .Y([1252]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10900 (.A([1250]), .B([1252]), .Y([1253]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10901 (.A([1254]), .B([1239]), .X([1255]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10902 (.A([496]), .B([1242]), .X([1256]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10903 (.A([1255]), .B([1256]), .Y([1257]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10904 (.A([1253]), .B([1257]), .X([1258]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10905 (.A([1259]), .B([1258]), .Y([1260]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10906 (.A([1248]), .B([1260]), .Y([1261]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10907 (.A([1262]), .B([1261]), .Y([1263]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10908 (.A([1264]), .B([1265]), .X([1266]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10909 (.A([1266]), .Y([1267]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10910 (.A([622]), .B([667]), .Y([1268]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10911 (.A([633]), .B([1268]), .X([1269]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10912 (.A([1186]), .B([1269]), .X([1270]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10913 (.A([1266]), .B([1270]), .X([1271]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10914 (.A([1196]), .B([1183]), .Y([1272]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10915 (.A([1272]), .Y([1273]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10916 (.A([1274]), .B([150]), .Y([1275]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10917 (.A([1276]), .B([1275]), .X([1277]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10918 (.A([662]), .B([693]), .Y([1278]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10919 (.A([1127]), .B([1278]), .X([1279]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10920 (.A([1277]), .B([1279]), .X([1280]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10921 (.A([1280]), .Y([1281]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10922 (.A([1263]), .B([1281]), .Y([1282]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10923 (.A([1271]), .B([1282]), .X([1283]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10924 (.A([1273]), .B([1283]), .X([1284]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10925 (.A([1284]), .Y([1285]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10926 (.A([1227]), .B([1285]), .Y([1286]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10927 (.A([1172]), .B([1286]), .X([1287]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10928 (.A([1288]), .B([1173]), .X([1289]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10929 (.A([1287]), .B([1289]), .Y([1290]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10930 (.A([1290]), .Y([1291]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10931 (.A([1178]), .B([1222]), .X([1292]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10932 (.A([1093]), .B([1292]), .X([1293]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10933 (.A([472]), .B([1293]), .Y([1294]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10934 (.A([172]), .B([1295]), .Y([1296]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10935 (.A([625]), .B([1296]), .X([1297]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10936 (.A([645]), .B([1157]), .X([1298]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10937 (.A([630]), .B([1127]), .X([1299]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10938 (.A([1298]), .B([1299]), .X([1300]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10939 (.A([1297]), .B([1300]), .X([1301]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10940 (.A([1132]), .B([1302]), .Y([1303]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10941 (.A([694]), .B([662]), .Y([1304]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10942 (.A([1304]), .Y([1305]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10943 (.A([1131]), .B([1304]), .X([1306]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10944 (.A([1303]), .B([1306]), .X([1307]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10945 (.A([1117]), .B([1307]), .X([1308]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10946 (.A([1301]), .B([1308]), .X([1309]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10947 (.A([562]), .B([1183]), .Y([1310]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10948 (.A([1122]), .B([1310]), .Y([1311]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10949 (.A([1311]), .Y([1312]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10950 (.A([1294]), .B([1312]), .Y([1313]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10951 (.A([1309]), .B([1313]), .X([1314]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10952 (.A([1173]), .B([1314]), .Y([1315]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10953 (.A([1316]), .B([1172]), .Y([1317]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10954 (.A([1315]), .B([1317]), .Y([1318]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10955 (.A([1053]), .B([1105]), .Y([1319]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10956 (.A([1102]), .B([1223]), .Y([1320]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10957 (.A([1319]), .B([1320]), .X([1321]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10958 (.A([1177]), .B([1321]), .X([1322]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10959 (.A([472]), .B([1322]), .Y([1323]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10960 (.A([644]), .B([1194]), .X([1324]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10961 (.A([1324]), .Y([1325]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10962 (.A([1198]), .B([1305]), .Y([1326]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10963 (.A([1325]), .B([1326]), .X([1327]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10964 (.A([1117]), .B([1327]), .X([1328]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10965 (.A([1130]), .B([469]), .Y([1329]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10966 (.A([1329]), .Y([1330]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10967 (.A([1331]), .B([1330]), .Y([1332]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10968 (.A([630]), .B([1149]), .X([1333]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10969 (.A([1332]), .B([1333]), .X([1334]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10970 (.A([1335]), .B([1155]), .X([1336]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10971 (.A([1190]), .B([1336]), .X([1337]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10972 (.A([1334]), .B([1337]), .X([1338]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10973 (.A([1328]), .B([1338]), .X([1339]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10974 (.A([1295]), .B([1261]), .X([1340]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10975 (.A([1312]), .B([1340]), .Y([1341]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10976 (.A([1339]), .B([1341]), .X([1342]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10977 (.A([1342]), .Y([1343]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10978 (.A([1323]), .B([1343]), .Y([1344]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10979 (.A([1173]), .B([1344]), .Y([1345]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10980 (.A([1346]), .B([1172]), .Y([1347]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10981 (.A([1345]), .B([1347]), .Y([1348]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10982 (.A([1349]), .B([1063]), .X([1350]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10983 (.A([1171]), .B([1350]), .Y([1351]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10984 (.A([1054]), .B([1351]), .X([1352]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10985 (.A([1220]), .B([1352]), .X([1353]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10986 (.A([472]), .B([1353]), .Y([1354]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10987 (.A([644]), .B([1195]), .X([1355]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10988 (.A([694]), .B([607]), .Y([1356]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10989 (.A([624]), .B([1156]), .Y([1357]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10990 (.A([1356]), .B([1357]), .X([1358]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10991 (.A([1359]), .B([1127]), .X([1360]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10992 (.A([1358]), .B([1360]), .X([1361]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10993 (.A([1336]), .B([1361]), .X([1362]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10994 (.A([1124]), .B([1355]), .Y([1363]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10995 (.A([1363]), .Y([1364]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10996 (.A([1354]), .B([1364]), .Y([1365]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10997 (.A([1362]), .B([1365]), .X([1366]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10998 (.A([1173]), .B([1366]), .Y([1367]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10999 (.A([1368]), .B([1172]), .Y([1369]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11000 (.A([1367]), .B([1369]), .Y([1370]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11001 (.A([1063]), .B([1170]), .Y([1371]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11002 (.A([1086]), .B([1179]), .X([1372]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11003 (.A([1371]), .B([1372]), .X([1373]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11004 (.A([472]), .B([1373]), .Y([1374]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11005 (.A([1134]), .B([1189]), .X([1375]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11006 (.A([697]), .B([1278]), .X([1376]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11007 (.A([1273]), .B([1376]), .X([1377]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11008 (.A([1375]), .B([1377]), .X([1378]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11009 (.A([1378]), .Y([1379]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11010 (.A([1374]), .B([1379]), .Y([1380]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11011 (.A([1140]), .B([1380]), .X([1381]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11012 (.A([1173]), .B([1381]), .Y([1382]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11013 (.A([1383]), .B([1172]), .Y([1384]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11014 (.A([1382]), .B([1384]), .Y([1385]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11015 (.A([1386]), .B([1387]), .X([1388]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11016 (.A([1047]), .B([1389]), .X([1390]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11017 (.A([1349]), .B([1069]), .X([1391]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11018 (.A([1391]), .Y([1392]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11019 (.A([1049]), .B([1393]), .X([1394]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11020 (.A([1395]), .B([1394]), .X([1396]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11021 (.A([1072]), .B([1397]), .X([1398]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11022 (.A([1055]), .B([1397]), .X([1399]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11023 (.A([1392]), .B([1399]), .X([1400]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11024 (.A([1390]), .B([1400]), .Y([1401]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11025 (.A([1396]), .B([1398]), .Y([1402]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11026 (.A([1401]), .B([1402]), .X([1403]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11027 (.A([1404]), .B([1403]), .X([1405]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11028 (.A([1406]), .B([1405]), .X([1407]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11029 (.A([1388]), .B([1407]), .Y([1408]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11030 (.A([1408]), .Y([1409]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11031 (.A([1410]), .B([1387]), .X([1411]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11032 (.A([1412]), .B([1413]), .X([1414]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11033 (.A([1085]), .B([1414]), .X([1415]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11034 (.A([1415]), .Y([1416]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11035 (.A([1078]), .B([1401]), .X([1417]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11036 (.A([1416]), .B([1417]), .X([1418]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11037 (.A([1404]), .B([1418]), .X([1419]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11038 (.A([1411]), .B([1419]), .Y([1420]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11039 (.A([1420]), .Y([1421]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11040 (.A([1422]), .B([1404]), .Y([1423]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11041 (.A([1395]), .B([1414]), .X([1424]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11042 (.A([1061]), .B([440]), .X([1425]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11043 (.A([1413]), .B([1425]), .X([1426]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11044 (.A([1426]), .Y([1427]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11045 (.A([1428]), .B([1424]), .Y([1429]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11046 (.A([1427]), .B([1429]), .X([1430]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11047 (.A([1431]), .B([1430]), .Y([1432]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11048 (.A([1387]), .B([1390]), .Y([1433]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11049 (.A([1433]), .Y([1434]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11050 (.A([1432]), .B([1434]), .Y([1435]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11051 (.A([1436]), .B([1425]), .Y([1437]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11052 (.A([1438]), .B([1437]), .Y([1439]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11053 (.A([1394]), .B([1439]), .Y([1440]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11054 (.A([1406]), .B([1440]), .X([1441]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11055 (.A([1435]), .B([1441]), .X([1442]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11056 (.A([1423]), .B([1442]), .Y([1443]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11057 (.A([1443]), .Y([1444]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11058 (.A([1085]), .B([1445]), .X([1446]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11059 (.A([1446]), .Y([1447]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11060 (.A([1435]), .B([1447]), .X([1448]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11061 (.A([1449]), .B([1387]), .X([1450]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11062 (.A([1448]), .B([1450]), .Y([1451]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11063 (.A([1451]), .Y([1452]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11064 (.A([1453]), .B([1387]), .X([1454]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11065 (.A([1455]), .B([1456]), .Y([1457]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11066 (.A([1073]), .B([1457]), .X([1458]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11067 (.A([1458]), .Y([1459]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11068 (.A([1460]), .B([1072]), .X([1461]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11069 (.A([1461]), .Y([1462]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11070 (.A([1463]), .B([1464]), .Y([1465]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11071 (.A([1462]), .B([1465]), .X([1466]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11072 (.A([1404]), .B([1466]), .X([1467]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11073 (.A([1459]), .B([1465]), .X([1468]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11074 (.A([1468]), .Y([1469]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11075 (.A([1459]), .B([1467]), .X([1470]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11076 (.A([1454]), .B([1470]), .Y([1471]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11077 (.A([1471]), .Y([1472]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11078 (.A([440]), .B([1473]), .X([1474]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11079 (.A([1474]), .Y([1475]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11080 (.A([445]), .B([1390]), .X([1476]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11081 (.A([1477]), .B([1073]), .X([1478]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11082 (.A([1479]), .B([1478]), .Y([1480]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11083 (.A([1480]), .Y([1481]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11084 (.A([1476]), .B([1481]), .Y([1482]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11085 (.A([1475]), .B([1482]), .X([1483]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11086 (.A([1484]), .B([1483]), .X([1485]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11087 (.A([1468]), .B([1485]), .X([1486]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11088 (.A([1387]), .B([1486]), .Y([1487]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11089 (.A([1488]), .B([1404]), .Y([1489]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11090 (.A([1487]), .B([1489]), .Y([1490]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11091 (.A([1491]), .B([1387]), .X([1492]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11092 (.A([1462]), .B([1486]), .X([1493]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11093 (.A([1387]), .B([1493]), .Y([1494]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11094 (.A([1072]), .B([1495]), .Y([1496]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11095 (.A([1497]), .B([1496]), .Y([1498]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11096 (.A([1498]), .Y([1499]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11097 (.A([1485]), .B([1499]), .X([1500]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11098 (.A([1494]), .B([1500]), .X([1501]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11099 (.A([1492]), .B([1501]), .Y([1502]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11100 (.A([1502]), .Y([1503]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11101 (.A([1504]), .B([1387]), .X([1505]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11102 (.A([1506]), .B([1458]), .X([1507]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11103 (.A([1507]), .Y([1508]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11104 (.A([1467]), .B([1508]), .X([1509]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11105 (.A([1469]), .B([1509]), .X([1510]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11106 (.A([1505]), .B([1510]), .Y([1511]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11107 (.A([1511]), .Y([1512]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11108 (.A([433]), .B([1513]), .Y([1514]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11109 (.A([148]), .B([645]), .X([1515]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11110 (.A([1066]), .B([647]), .Y([1516]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11111 (.A([1517]), .B([663]), .X([1518]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11112 (.A([456]), .B([1518]), .X([1519]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11113 (.A([1516]), .B([1519]), .X([1520]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11114 (.A([1515]), .B([1520]), .X([1521]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11115 (.A([1521]), .Y([1522]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11116 (.A([1523]), .B([577]), .Y([1524]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11117 (.A([539]), .B([1525]), .X([1526]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11118 (.A([44]), .B([1526]), .Y([1527]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11119 (.A([1243]), .B([1526]), .X([1528]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11120 (.A([1527]), .B([1528]), .Y([1529]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11121 (.A([544]), .B([1529]), .X([1530]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11122 (.A([1531]), .B([544]), .Y([1532]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11123 (.A([1530]), .B([1532]), .Y([1533]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11124 (.A([1523]), .B([1533]), .X([1534]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11125 (.A([1524]), .B([1534]), .Y([1535]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11126 (.A([1517]), .B([1535]), .Y([1536]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11127 (.A([1536]), .Y([1537]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11128 (.A([550]), .B([1515]), .Y([1538]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11129 (.A([1538]), .Y([1539]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11130 (.A([607]), .B([667]), .Y([1540]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11131 (.A([628]), .B([1540]), .X([1541]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11132 (.A([1139]), .B([1541]), .X([1542]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11133 (.A([539]), .B([1543]), .X([1544]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11134 (.A([539]), .B([456]), .Y([1545]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11135 (.A([1544]), .B([1545]), .Y([1546]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11136 (.A([1523]), .B([1546]), .X([1547]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11137 (.A([1524]), .B([1547]), .Y([1548]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11138 (.A([663]), .B([1548]), .Y([1549]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11139 (.A([1267]), .B([1549]), .Y([1550]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11140 (.A([1542]), .B([1550]), .X([1551]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11141 (.A([1539]), .B([1551]), .X([1552]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11142 (.A([1537]), .B([1552]), .X([1553]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11143 (.A([1522]), .B([1553]), .X([1554]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11144 (.A([1555]), .B([1518]), .Y([1556]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11145 (.A([1519]), .B([1556]), .Y([1557]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11146 (.A([1557]), .Y([1558]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11147 (.A([1554]), .B([1558]), .X([1559]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11148 (.A([1274]), .B([1161]), .Y([1560]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11149 (.A([661]), .B([1560]), .X([1561]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11150 (.A([695]), .B([1561]), .X([1562]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11151 (.A([1563]), .B([1303]), .X([1564]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11152 (.A([1565]), .B([1564]), .X([1566]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11153 (.A([1562]), .B([1566]), .X([1567]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11154 (.A([1525]), .B([1113]), .X([1568]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11155 (.A([1568]), .Y([1569]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11156 (.A([1567]), .B([1569]), .X([1570]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11157 (.A([1570]), .Y([1571]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11158 (.A([894]), .B([1571]), .X([1572]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11159 (.A([607]), .B([632]), .Y([1573]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11160 (.A([628]), .B([1573]), .X([1574]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11161 (.A([626]), .B([1574]), .X([1575]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11162 (.A([1517]), .B([1516]), .X([1576]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11163 (.A([1295]), .B([662]), .Y([1577]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11164 (.A([1578]), .B([1577]), .X([1579]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11165 (.A([1576]), .B([1579]), .X([1580]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11166 (.A([1575]), .B([1580]), .X([1581]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11167 (.A([1567]), .B([1581]), .X([1582]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11168 (.A([1582]), .Y([1583]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11169 (.A([1525]), .B([44]), .Y([1584]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11170 (.A([1113]), .B([1584]), .X([1585]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11171 (.A([1582]), .B([1585]), .Y([1586]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11172 (.A([234]), .B([1575]), .Y([1587]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11173 (.A([419]), .B([1577]), .Y([1588]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11174 (.A([424]), .B([1588]), .Y([1589]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11175 (.A([1589]), .Y([1590]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11176 (.A([1587]), .B([1590]), .Y([1591]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11177 (.A([1586]), .B([1591]), .X([1592]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11178 (.A([1592]), .Y([1593]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11179 (.A([1572]), .B([1593]), .Y([1594]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11180 (.A([1504]), .B([1518]), .Y([1595]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11181 (.A([1595]), .Y([1596]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11182 (.A([1491]), .B([1518]), .Y([1597]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11183 (.A([1597]), .Y([1598]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11184 (.A([1599]), .B([1187]), .X([1600]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11185 (.A([1149]), .B([1600]), .X([1601]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11186 (.A([148]), .B([1601]), .X([1602]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11187 (.A([1531]), .B([663]), .X([1603]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11188 (.A([1576]), .B([1603]), .X([1604]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11189 (.A([1604]), .Y([1605]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11190 (.A([1602]), .B([1605]), .X([1606]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11191 (.A([1598]), .B([1606]), .X([1607]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11192 (.A([1596]), .B([1606]), .X([1608]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11193 (.A([1596]), .B([1607]), .X([1609]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11194 (.A([627]), .B([662]), .Y([1610]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11195 (.A([620]), .B([1610]), .X([1611]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11196 (.A([1516]), .B([1573]), .X([1612]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11197 (.A([1611]), .B([1612]), .X([1613]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11198 (.A([1297]), .B([1564]), .X([1614]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11199 (.A([1613]), .B([1614]), .X([1615]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11200 (.A([1562]), .B([1615]), .X([1616]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11201 (.A([1616]), .Y([1617]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11202 (.A([419]), .B([1617]), .Y([1618]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11203 (.A([232]), .B([1262]), .Y([1619]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11204 (.A([1618]), .B([1619]), .Y([1620]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11205 (.A([1620]), .Y([1621]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11206 (.A([1608]), .B([1621]), .X([1622]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11207 (.A([1607]), .B([1620]), .X([1623]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11208 (.A([1622]), .B([1623]), .Y([1624]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11209 (.A([1609]), .B([1624]), .Y([1625]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11210 (.A([1594]), .B([1622]), .X([1626]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11211 (.A([1626]), .Y([1627]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11212 (.A([1594]), .B([1625]), .Y([1628]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11213 (.A([1558]), .B([1628]), .Y([1629]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11214 (.A([1627]), .B([1629]), .X([1630]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11215 (.A([1559]), .B([1630]), .Y([1631]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11216 (.A([1520]), .B([1602]), .X([1632]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11217 (.A([1453]), .B([1518]), .Y([1633]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11218 (.A([1632]), .B([1633]), .Y([1634]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11219 (.A([583]), .B([148]), .Y([1635]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11220 (.A([1488]), .B([1518]), .Y([1636]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11221 (.A([1635]), .B([1636]), .Y([1637]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11222 (.A([1601]), .B([1637]), .X([1638]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11223 (.A([1638]), .Y([1639]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11224 (.A([1632]), .B([1639]), .Y([1640]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11225 (.A([1634]), .B([1638]), .X([1641]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11226 (.A([1620]), .B([1641]), .Y([1642]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11227 (.A([1634]), .B([1639]), .X([1643]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11228 (.A([1621]), .B([1643]), .Y([1644]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11229 (.A([1642]), .B([1644]), .Y([1645]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11230 (.A([1631]), .B([1645]), .Y([1646]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11231 (.A([1633]), .B([1640]), .X([1647]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11232 (.A([1647]), .Y([1648]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11233 (.A([1645]), .B([1647]), .Y([1649]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11234 (.A([1649]), .Y([1650]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11235 (.A([1646]), .B([1649]), .Y([1651]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11236 (.A([433]), .B([1651]), .X([1652]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11237 (.A([1514]), .B([1652]), .Y([1653]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11238 (.A([39]), .B([234]), .X([1654]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11239 (.A([1033]), .B([1616]), .X([1655]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11240 (.A([211]), .B([1262]), .Y([1656]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11241 (.A([1655]), .B([1656]), .Y([1657]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11242 (.A([1657]), .Y([1658]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11243 (.A([1643]), .B([1657]), .X([1659]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11244 (.A([1641]), .B([1658]), .X([1660]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11245 (.A([1659]), .B([1660]), .Y([1661]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11246 (.A([1648]), .B([1661]), .X([1662]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11247 (.A([865]), .B([1571]), .X([1663]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11248 (.A([213]), .B([1575]), .Y([1664]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11249 (.A([398]), .B([1577]), .Y([1665]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11250 (.A([401]), .B([1665]), .Y([1666]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11251 (.A([1585]), .B([1664]), .Y([1667]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11252 (.A([1583]), .B([1667]), .X([1668]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11253 (.A([1666]), .B([1668]), .X([1669]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11254 (.A([1669]), .Y([1670]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11255 (.A([1663]), .B([1670]), .Y([1671]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11256 (.A([1671]), .Y([1672]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11257 (.A([1608]), .B([1658]), .X([1673]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11258 (.A([1672]), .B([1673]), .Y([1674]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11259 (.A([1674]), .Y([1675]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11260 (.A([1607]), .B([1657]), .X([1676]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11261 (.A([1673]), .B([1676]), .Y([1677]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11262 (.A([1609]), .B([1677]), .Y([1678]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11263 (.A([1672]), .B([1678]), .X([1679]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11264 (.A([1557]), .B([1594]), .Y([1680]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11265 (.A([1558]), .B([1679]), .Y([1681]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11266 (.A([1675]), .B([1681]), .X([1682]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11267 (.A([1680]), .B([1682]), .Y([1683]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11268 (.A([1662]), .B([1683]), .Y([1684]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11269 (.A([1028]), .B([1616]), .X([1685]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11270 (.A([189]), .B([1262]), .Y([1686]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11271 (.A([1685]), .B([1686]), .Y([1687]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11272 (.A([1687]), .Y([1688]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11273 (.A([1641]), .B([1687]), .Y([1689]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11274 (.A([1643]), .B([1688]), .Y([1690]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11275 (.A([1689]), .B([1690]), .Y([1691]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11276 (.A([1647]), .B([1691]), .Y([1692]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11277 (.A([1692]), .Y([1693]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11278 (.A([836]), .B([1571]), .X([1694]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11279 (.A([191]), .B([1575]), .Y([1695]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11280 (.A([375]), .B([1577]), .Y([1696]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11281 (.A([380]), .B([1696]), .Y([1697]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11282 (.A([1697]), .Y([1698]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11283 (.A([1695]), .B([1698]), .Y([1699]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11284 (.A([1586]), .B([1699]), .X([1700]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11285 (.A([1700]), .Y([1701]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11286 (.A([1694]), .B([1701]), .Y([1702]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11287 (.A([1608]), .B([1688]), .X([1703]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11288 (.A([1607]), .B([1687]), .X([1704]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11289 (.A([1703]), .B([1704]), .Y([1705]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11290 (.A([1609]), .B([1705]), .Y([1706]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11291 (.A([1702]), .B([1703]), .X([1707]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11292 (.A([1702]), .B([1706]), .Y([1708]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11293 (.A([1707]), .B([1708]), .Y([1709]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11294 (.A([1557]), .B([1709]), .X([1710]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11295 (.A([1558]), .B([1671]), .X([1711]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11296 (.A([1710]), .B([1711]), .Y([1712]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11297 (.A([1693]), .B([1712]), .X([1713]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11298 (.A([352]), .B([1617]), .Y([1714]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11299 (.A([167]), .B([1262]), .Y([1715]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11300 (.A([1714]), .B([1715]), .Y([1716]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11301 (.A([1716]), .Y([1717]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11302 (.A([1643]), .B([1716]), .X([1718]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11303 (.A([1641]), .B([1717]), .X([1719]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11304 (.A([1718]), .B([1719]), .Y([1720]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11305 (.A([1648]), .B([1720]), .X([1721]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11306 (.A([807]), .B([1571]), .X([1722]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11307 (.A([169]), .B([1575]), .Y([1723]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11308 (.A([352]), .B([1577]), .Y([1724]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11309 (.A([358]), .B([1724]), .Y([1725]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11310 (.A([1725]), .Y([1726]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11311 (.A([1723]), .B([1726]), .Y([1727]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11312 (.A([1586]), .B([1727]), .X([1728]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11313 (.A([1728]), .Y([1729]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11314 (.A([1722]), .B([1729]), .Y([1730]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11315 (.A([1608]), .B([1717]), .X([1731]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11316 (.A([1731]), .Y([1732]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11317 (.A([1607]), .B([1716]), .X([1733]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11318 (.A([1731]), .B([1733]), .Y([1734]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11319 (.A([1609]), .B([1734]), .Y([1735]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11320 (.A([1735]), .Y([1736]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11321 (.A([1730]), .B([1736]), .Y([1737]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11322 (.A([1730]), .B([1732]), .X([1738]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11323 (.A([1738]), .Y([1739]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11324 (.A([1557]), .B([1702]), .Y([1740]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11325 (.A([1558]), .B([1737]), .Y([1741]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11326 (.A([1739]), .B([1741]), .X([1742]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11327 (.A([1740]), .B([1742]), .Y([1743]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11328 (.A([1721]), .B([1743]), .Y([1744]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11329 (.A([468]), .B([1616]), .X([1745]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11330 (.A([142]), .B([1262]), .Y([1746]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11331 (.A([1745]), .B([1746]), .Y([1747]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11332 (.A([1747]), .Y([1748]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11333 (.A([1641]), .B([1747]), .Y([1749]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11334 (.A([1643]), .B([1748]), .Y([1750]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11335 (.A([1749]), .B([1750]), .Y([1751]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11336 (.A([1647]), .B([1751]), .Y([1752]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11337 (.A([1752]), .Y([1753]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11338 (.A([778]), .B([1571]), .X([1754]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11339 (.A([145]), .B([1575]), .Y([1755]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11340 (.A([329]), .B([1577]), .Y([1756]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11341 (.A([334]), .B([1756]), .Y([1757]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11342 (.A([1757]), .Y([1758]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11343 (.A([1755]), .B([1758]), .Y([1759]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11344 (.A([1586]), .B([1759]), .X([1760]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11345 (.A([1760]), .Y([1761]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11346 (.A([1754]), .B([1761]), .Y([1762]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11347 (.A([1608]), .B([1748]), .X([1763]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11348 (.A([1607]), .B([1747]), .X([1764]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11349 (.A([1763]), .B([1764]), .Y([1765]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11350 (.A([1609]), .B([1765]), .Y([1766]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11351 (.A([1762]), .B([1763]), .X([1767]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11352 (.A([1762]), .B([1766]), .Y([1768]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11353 (.A([1767]), .B([1768]), .Y([1769]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11354 (.A([1557]), .B([1769]), .X([1770]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11355 (.A([1558]), .B([1730]), .X([1771]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11356 (.A([1770]), .B([1771]), .Y([1772]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11357 (.A([1753]), .B([1772]), .X([1773]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11358 (.A([1751]), .B([1772]), .Y([1774]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11359 (.A([1773]), .B([1774]), .Y([1775]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11360 (.A([1775]), .Y([1776]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11361 (.A([1015]), .B([1616]), .X([1777]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11362 (.A([138]), .B([1262]), .Y([1778]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11363 (.A([1777]), .B([1778]), .Y([1779]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11364 (.A([1779]), .Y([1780]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11365 (.A([1641]), .B([1779]), .Y([1781]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11366 (.A([1643]), .B([1780]), .Y([1782]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11367 (.A([1781]), .B([1782]), .Y([1783]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11368 (.A([1647]), .B([1783]), .Y([1784]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11369 (.A([1784]), .Y([1785]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11370 (.A([749]), .B([1571]), .X([1786]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11371 (.A([518]), .B([1575]), .Y([1787]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11372 (.A([305]), .B([1577]), .Y([1788]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11373 (.A([1585]), .B([1788]), .Y([1789]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11374 (.A([312]), .B([1789]), .X([1790]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11375 (.A([1790]), .Y([1791]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11376 (.A([1787]), .B([1791]), .Y([1792]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11377 (.A([1583]), .B([1792]), .X([1793]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11378 (.A([1793]), .Y([1794]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11379 (.A([1786]), .B([1794]), .Y([1795]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11380 (.A([1608]), .B([1780]), .X([1796]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11381 (.A([1607]), .B([1779]), .X([1797]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11382 (.A([1796]), .B([1797]), .Y([1798]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11383 (.A([1609]), .B([1798]), .Y([1799]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11384 (.A([1795]), .B([1796]), .X([1800]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11385 (.A([1795]), .B([1799]), .Y([1801]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11386 (.A([1800]), .B([1801]), .Y([1802]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11387 (.A([1557]), .B([1802]), .X([1803]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11388 (.A([1558]), .B([1762]), .X([1804]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11389 (.A([1803]), .B([1804]), .Y([1805]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11390 (.A([1785]), .B([1805]), .X([1806]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11391 (.A([508]), .B([1616]), .X([1807]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11392 (.A([721]), .B([1262]), .Y([1808]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11393 (.A([1807]), .B([1808]), .Y([1809]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11394 (.A([1809]), .Y([1810]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11395 (.A([1643]), .B([1809]), .X([1811]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11396 (.A([1641]), .B([1810]), .X([1812]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11397 (.A([1811]), .B([1812]), .Y([1813]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11398 (.A([1648]), .B([1813]), .X([1814]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11399 (.A([718]), .B([1571]), .X([1815]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11400 (.A([286]), .B([1575]), .Y([1816]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11401 (.A([281]), .B([1577]), .Y([1817]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11402 (.A([285]), .B([1582]), .Y([1818]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11403 (.A([1585]), .B([1817]), .Y([1819]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11404 (.A([1819]), .Y([1820]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11405 (.A([1816]), .B([1820]), .Y([1821]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11406 (.A([1818]), .B([1821]), .X([1822]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11407 (.A([1822]), .Y([1823]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11408 (.A([1815]), .B([1823]), .Y([1824]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11409 (.A([1608]), .B([1810]), .X([1825]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11410 (.A([1607]), .B([1809]), .X([1826]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11411 (.A([1825]), .B([1826]), .Y([1827]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11412 (.A([1609]), .B([1827]), .Y([1828]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11413 (.A([1824]), .B([1828]), .Y([1829]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11414 (.A([1824]), .B([1825]), .X([1830]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11415 (.A([1829]), .B([1830]), .Y([1831]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11416 (.A([1558]), .B([1831]), .Y([1832]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11417 (.A([1557]), .B([1795]), .Y([1833]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11418 (.A([1832]), .B([1833]), .Y([1834]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11419 (.A([1814]), .B([1834]), .Y([1835]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11420 (.A([567]), .B([1616]), .X([1836]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11421 (.A([675]), .B([1262]), .Y([1837]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11422 (.A([1836]), .B([1837]), .Y([1838]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11423 (.A([1838]), .Y([1839]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11424 (.A([1643]), .B([1838]), .X([1840]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11425 (.A([1641]), .B([1839]), .X([1841]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11426 (.A([1840]), .B([1841]), .Y([1842]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11427 (.A([1648]), .B([1842]), .X([1843]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11428 (.A([1557]), .B([1824]), .Y([1844]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11429 (.A([602]), .B([1570]), .Y([1845]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11430 (.A([516]), .B([1575]), .Y([1846]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11431 (.A([256]), .B([1577]), .Y([1847]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11432 (.A([260]), .B([1847]), .Y([1848]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11433 (.A([1848]), .Y([1849]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11434 (.A([1846]), .B([1849]), .Y([1850]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11435 (.A([1586]), .B([1850]), .X([1851]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11436 (.A([1851]), .Y([1852]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11437 (.A([1845]), .B([1852]), .Y([1853]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11438 (.A([1608]), .B([1839]), .X([1854]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11439 (.A([1607]), .B([1838]), .X([1855]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11440 (.A([1854]), .B([1855]), .Y([1856]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11441 (.A([1609]), .B([1856]), .Y([1857]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11442 (.A([1853]), .B([1854]), .X([1858]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11443 (.A([1853]), .B([1857]), .Y([1859]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11444 (.A([1858]), .B([1859]), .Y([1860]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11445 (.A([1558]), .B([1860]), .Y([1861]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11446 (.A([1844]), .B([1861]), .Y([1862]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11447 (.A([1843]), .B([1862]), .Y([1863]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11448 (.A([1842]), .B([1862]), .X([1864]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11449 (.A([1863]), .B([1864]), .Y([1865]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11450 (.A([1634]), .B([1640]), .Y([1866]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11451 (.A([1558]), .B([1866]), .Y([1867]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11452 (.A([1554]), .B([1867]), .X([1868]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11453 (.A([456]), .B([1867]), .Y([1869]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11454 (.A([1868]), .B([1869]), .Y([1870]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11455 (.A([1865]), .B([1870]), .X([1871]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11456 (.A([1863]), .B([1871]), .Y([1872]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11457 (.A([1813]), .B([1834]), .X([1873]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11458 (.A([1835]), .B([1873]), .Y([1874]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11459 (.A([1874]), .Y([1875]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11460 (.A([1872]), .B([1875]), .Y([1876]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11461 (.A([1835]), .B([1876]), .Y([1877]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11462 (.A([1783]), .B([1805]), .Y([1878]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11463 (.A([1806]), .B([1878]), .Y([1879]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11464 (.A([1879]), .Y([1880]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11465 (.A([1877]), .B([1880]), .Y([1881]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11466 (.A([1806]), .B([1881]), .Y([1882]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11467 (.A([1776]), .B([1882]), .Y([1883]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11468 (.A([1776]), .B([1882]), .X([1884]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11469 (.A([1883]), .B([1884]), .Y([1885]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11470 (.A([1886]), .B([1517]), .Y([1887]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11471 (.A([1887]), .Y([1888]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11472 (.A([1877]), .B([1880]), .X([1889]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11473 (.A([1881]), .B([1889]), .Y([1890]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11474 (.A([1872]), .B([1875]), .X([1891]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11475 (.A([1876]), .B([1891]), .Y([1892]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11476 (.A([1890]), .B([1892]), .Y([1893]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11477 (.A([1888]), .B([1893]), .Y([1894]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11478 (.A([1885]), .B([1894]), .X([1895]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11479 (.A([1773]), .B([1883]), .Y([1896]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11480 (.A([1896]), .Y([1897]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11481 (.A([1895]), .B([1897]), .Y([1898]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11482 (.A([1720]), .B([1743]), .X([1899]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11483 (.A([1744]), .B([1899]), .Y([1900]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11484 (.A([1900]), .Y([1901]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11485 (.A([1898]), .B([1901]), .Y([1902]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11486 (.A([1744]), .B([1902]), .Y([1903]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11487 (.A([1691]), .B([1712]), .Y([1904]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11488 (.A([1713]), .B([1904]), .Y([1905]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11489 (.A([1905]), .Y([1906]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11490 (.A([1903]), .B([1906]), .Y([1907]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11491 (.A([1713]), .B([1907]), .Y([1908]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11492 (.A([1661]), .B([1683]), .X([1909]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11493 (.A([1684]), .B([1909]), .Y([1910]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11494 (.A([1910]), .Y([1911]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11495 (.A([1908]), .B([1911]), .Y([1912]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11496 (.A([1684]), .B([1912]), .Y([1913]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11497 (.A([1631]), .B([1650]), .X([1914]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11498 (.A([1914]), .Y([1915]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11499 (.A([1646]), .B([1914]), .Y([1916]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11500 (.A([1913]), .B([1916]), .Y([1917]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11501 (.A([1913]), .B([1916]), .X([1918]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11502 (.A([1917]), .B([1918]), .Y([1919]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11503 (.A([433]), .B([1919]), .X([1920]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11504 (.A([1654]), .B([1920]), .Y([1921]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11505 (.A([1921]), .Y([1922]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11506 (.A([433]), .B([1923]), .Y([1924]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11507 (.A([39]), .B([1898]), .Y([1925]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11508 (.A([1924]), .B([1925]), .Y([1926]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11509 (.A([1865]), .B([1870]), .Y([1927]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11510 (.A([1871]), .B([1927]), .Y([1928]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11511 (.A([39]), .B([1928]), .Y([1929]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11512 (.A([39]), .B([516]), .X([1930]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11513 (.A([1929]), .B([1930]), .Y([1931]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11514 (.A([1931]), .Y([1932]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11515 (.A([39]), .B([286]), .X([1933]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11516 (.A([39]), .B([1892]), .Y([1934]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11517 (.A([1933]), .B([1934]), .Y([1935]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11518 (.A([1935]), .Y([1936]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11519 (.A([39]), .B([518]), .X([1937]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11520 (.A([39]), .B([1890]), .Y([1938]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11521 (.A([1937]), .B([1938]), .Y([1939]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11522 (.A([1939]), .Y([1940]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11523 (.A([39]), .B([145]), .X([1941]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11524 (.A([39]), .B([1885]), .Y([1942]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11525 (.A([1941]), .B([1942]), .Y([1943]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11526 (.A([1943]), .Y([1944]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11527 (.A([1898]), .B([1901]), .X([1945]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11528 (.A([1902]), .B([1945]), .Y([1946]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11529 (.A([39]), .B([1946]), .Y([1947]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11530 (.A([39]), .B([169]), .X([1948]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11531 (.A([1947]), .B([1948]), .Y([1949]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11532 (.A([1949]), .Y([1950]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11533 (.A([1903]), .B([1906]), .X([1951]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11534 (.A([1907]), .B([1951]), .Y([1952]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11535 (.A([39]), .B([191]), .X([1953]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11536 (.A([39]), .B([1952]), .Y([1954]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11537 (.A([1953]), .B([1954]), .Y([1955]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11538 (.A([1955]), .Y([1956]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11539 (.A([1908]), .B([1911]), .X([1957]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11540 (.A([1912]), .B([1957]), .Y([1958]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11541 (.A([39]), .B([213]), .X([1959]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11542 (.A([39]), .B([1958]), .Y([1960]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11543 (.A([1959]), .B([1960]), .Y([1961]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11544 (.A([1961]), .Y([1962]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11545 (.A([433]), .B([1963]), .Y([1964]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11546 (.A([39]), .B([1594]), .Y([1965]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11547 (.A([1964]), .B([1965]), .Y([1966]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11548 (.A([39]), .B([550]), .X([1967]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11549 (.A([1558]), .B([1853]), .X([1968]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11550 (.A([456]), .B([1556]), .Y([1969]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11551 (.A([1968]), .B([1969]), .Y([1970]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11552 (.A([1913]), .B([1915]), .X([1971]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11553 (.A([1646]), .B([1971]), .Y([1972]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11554 (.A([1970]), .B([1972]), .X([1973]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11555 (.A([1970]), .B([1972]), .Y([1974]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11556 (.A([1973]), .B([1974]), .Y([1975]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11557 (.A([1952]), .B([1958]), .Y([1976]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11558 (.A([1888]), .B([1976]), .Y([1977]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11559 (.A([39]), .B([1977]), .Y([1978]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11560 (.A([1920]), .B([1978]), .Y([1979]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11561 (.A([1975]), .B([1979]), .Y([1980]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11562 (.A([1967]), .B([1980]), .Y([1981]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11563 (.A([1981]), .Y([1982]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11564 (.A([1983]), .B([1125]), .X([1984]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11565 (.A([38]), .B([1985]), .Y([1986]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11566 (.A([1531]), .B([1986]), .X([1987]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11567 (.A([1988]), .B([1986]), .Y([1989]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11568 (.A([1987]), .B([1989]), .Y([1990]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11569 (.A([1984]), .B([1990]), .Y([1991]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11570 (.A([1991]), .Y([1992]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11571 (.A([456]), .B([1066]), .X([1993]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11572 (.A([1993]), .Y([1994]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11573 (.A([1995]), .B([1066]), .Y([1996]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11574 (.A([3]), .B([1996]), .Y([1997]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11575 (.A([1994]), .B([1997]), .X([1998]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11576 (.A([1404]), .B([1001]), .Y([1999]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11577 (.A([2000]), .B([1999]), .X([2001]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11578 (.A([696]), .B([1993]), .Y([2002]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11579 (.A([1531]), .B([695]), .Y([2003]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11580 (.A([2002]), .B([2003]), .Y([2004]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11581 (.A([1999]), .B([2004]), .Y([2005]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11582 (.A([2001]), .B([2005]), .Y([2006]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11583 (.A([1002]), .B([2006]), .X([2007]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11584 (.A([2007]), .Y([2008]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11585 (.A([2009]), .B([476]), .Y([2010]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11586 (.A([309]), .B([476]), .X([2011]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11587 (.A([2010]), .B([2011]), .Y([2012]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11588 (.A([660]), .B([2012]), .Y([2013]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11589 (.A([60]), .B([2014]), .Y([2015]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11590 (.A([2016]), .B([2009]), .Y([2017]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11591 (.A([2015]), .B([2017]), .Y([2018]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11592 (.A([2019]), .B([2018]), .Y([2020]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11593 (.A([2021]), .B([44]), .Y([2022]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11594 (.A([2020]), .B([2022]), .Y([2023]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11595 (.A([661]), .B([2023]), .Y([2024]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11596 (.A([2013]), .B([2024]), .Y([2025]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11597 (.A([469]), .B([2025]), .Y([2026]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11598 (.A([1015]), .B([469]), .X([2027]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11599 (.A([1125]), .B([2027]), .Y([2028]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11600 (.A([2028]), .Y([2029]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11601 (.A([2026]), .B([2029]), .Y([2030]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11602 (.A([1118]), .B([1183]), .X([2031]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11603 (.A([1193]), .B([2031]), .Y([2032]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11604 (.A([491]), .B([1601]), .X([2033]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11605 (.A([2033]), .Y([2034]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11606 (.A([456]), .B([2031]), .X([2035]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11607 (.A([2032]), .B([2035]), .Y([2036]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11608 (.A([2033]), .B([2036]), .X([116]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11609 (.A([602]), .B([2034]), .Y([2037]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11610 (.A([2038]), .B([2039]), .X([2040]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11611 (.A([150]), .B([2040]), .Y([2041]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11612 (.A([577]), .B([2041]), .Y([2042]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11613 (.A([2043]), .B([2039]), .X([2044]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11614 (.A([490]), .B([2044]), .Y([2045]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11615 (.A([516]), .B([2045]), .Y([2046]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11616 (.A([1274]), .B([1160]), .Y([2047]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11617 (.A([253]), .B([2047]), .Y([2048]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11618 (.A([675]), .B([1149]), .Y([2049]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11619 (.A([2042]), .B([2049]), .Y([2050]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11620 (.A([2046]), .B([2048]), .Y([2051]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11621 (.A([2051]), .Y([2052]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11622 (.A([2037]), .B([2052]), .Y([2053]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11623 (.A([2050]), .B([2053]), .X([108]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11624 (.A([718]), .B([2033]), .X([2054]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11625 (.A([286]), .B([2045]), .Y([2055]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11626 (.A([2055]), .Y([2056]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11627 (.A([531]), .B([2041]), .Y([2057]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11628 (.A([279]), .B([2047]), .Y([2058]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11629 (.A([721]), .B([1149]), .Y([2059]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11630 (.A([2058]), .B([2059]), .Y([2060]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11631 (.A([2060]), .Y([2061]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11632 (.A([2057]), .B([2061]), .Y([2062]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11633 (.A([2056]), .B([2062]), .X([2063]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11634 (.A([2063]), .Y([2064]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11635 (.A([2054]), .B([2064]), .Y([109]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11636 (.A([749]), .B([2033]), .X([2065]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11637 (.A([2009]), .B([2041]), .Y([2066]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11638 (.A([2066]), .Y([2067]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11639 (.A([518]), .B([2045]), .Y([2068]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11640 (.A([138]), .B([1149]), .Y([2069]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11641 (.A([303]), .B([2047]), .Y([2070]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11642 (.A([2069]), .B([2070]), .Y([2071]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11643 (.A([2071]), .Y([2072]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11644 (.A([2068]), .B([2072]), .Y([2073]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11645 (.A([2067]), .B([2073]), .X([2074]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11646 (.A([2074]), .Y([2075]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11647 (.A([2065]), .B([2075]), .Y([110]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11648 (.A([778]), .B([2033]), .X([2076]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11649 (.A([145]), .B([2045]), .Y([2077]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11650 (.A([474]), .B([2041]), .Y([2078]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11651 (.A([327]), .B([2047]), .Y([2079]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11652 (.A([142]), .B([1149]), .Y([2080]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11653 (.A([2078]), .B([2080]), .Y([2081]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11654 (.A([2077]), .B([2079]), .Y([2082]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11655 (.A([2082]), .Y([2083]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11656 (.A([2076]), .B([2083]), .Y([2084]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11657 (.A([2081]), .B([2084]), .X([111]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11658 (.A([807]), .B([2033]), .X([2085]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11659 (.A([169]), .B([2045]), .Y([2086]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11660 (.A([2086]), .Y([2087]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11661 (.A([349]), .B([2047]), .Y([2088]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11662 (.A([167]), .B([1149]), .Y([2089]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11663 (.A([2088]), .B([2089]), .Y([2090]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11664 (.A([1531]), .B([2040]), .X([2091]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11665 (.A([2092]), .B([150]), .X([2093]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11666 (.A([2091]), .B([2093]), .Y([2094]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11667 (.A([2090]), .B([2094]), .X([2095]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11668 (.A([2087]), .B([2095]), .X([2096]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11669 (.A([2096]), .Y([2097]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11670 (.A([2085]), .B([2097]), .Y([112]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11671 (.A([836]), .B([2033]), .X([2098]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11672 (.A([191]), .B([2045]), .Y([2099]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11673 (.A([2099]), .Y([2100]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11674 (.A([150]), .B([2091]), .Y([2101]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11675 (.A([189]), .B([1149]), .Y([2102]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11676 (.A([373]), .B([2047]), .Y([2103]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11677 (.A([2102]), .B([2103]), .Y([2104]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11678 (.A([2101]), .B([2104]), .X([2105]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11679 (.A([2100]), .B([2105]), .X([2106]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11680 (.A([2106]), .Y([2107]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11681 (.A([2098]), .B([2107]), .Y([113]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11682 (.A([865]), .B([2033]), .X([2108]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11683 (.A([213]), .B([2045]), .Y([2109]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11684 (.A([2110]), .B([2041]), .Y([2111]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11685 (.A([2111]), .Y([2112]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11686 (.A([211]), .B([1149]), .Y([2113]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11687 (.A([2113]), .Y([2114]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11688 (.A([396]), .B([2047]), .Y([2115]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11689 (.A([2109]), .B([2115]), .Y([2116]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11690 (.A([2114]), .B([2116]), .X([2117]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11691 (.A([2112]), .B([2117]), .X([2118]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11692 (.A([2118]), .Y([2119]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11693 (.A([2108]), .B([2119]), .Y([114]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11694 (.A([894]), .B([2033]), .X([2120]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11695 (.A([2121]), .B([2041]), .Y([2122]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11696 (.A([2122]), .Y([2123]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11697 (.A([236]), .B([2044]), .X([2124]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11698 (.A([499]), .B([2124]), .Y([2125]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11699 (.A([417]), .B([2047]), .Y([2126]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11700 (.A([232]), .B([1149]), .Y([2127]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11701 (.A([2126]), .B([2127]), .Y([2128]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11702 (.A([2125]), .B([2128]), .X([2129]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11703 (.A([2123]), .B([2129]), .X([2130]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11704 (.A([2130]), .Y([2131]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11705 (.A([2120]), .B([2131]), .Y([115]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11706 (.A([546]), .B([474]), .Y([2132]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11707 (.A([2132]), .Y([2133]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9277 (.A([2134]), .Y([705]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9278 (.A([2135]), .Y([595]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9279 (.A([2136]), .Y([587]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9280 (.A([2110]), .Y([1254]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9281 (.A([1988]), .Y([1983]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9282 (.A([60]), .Y([1531]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9283 (.A([462]), .Y([2137]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9284 (.A([2043]), .Y([2038]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9285 (.A([453]), .Y([459]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9286 (.A([2021]), .Y([2019]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9287 (.A([2014]), .Y([2016]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9288 (.A([2138]), .Y([2139]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9289 (.A([544]), .Y([484]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9290 (.A([39]), .Y([433]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9291 (.A([448]), .Y([1259]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9292 (.A([2121]), .Y([496]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9293 (.A([531]), .Y([1240]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9294 (.A([577]), .Y([1243]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9295 (.A([1006]), .Y([2140]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9296 (.A([1010]), .Y([2141]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9297 (.A([1013]), .Y([2142]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9298 (.A([1019]), .Y([2143]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9299 (.A([1023]), .Y([2144]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9300 (.A([1031]), .Y([2145]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9301 (.A([1036]), .Y([2146]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9302 (.A([2147]), .Y([1422]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9303 (.A([234]), .Y([236]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9304 (.A([516]), .Y([263]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9305 (.A([518]), .Y([309]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9306 (.A([169]), .Y([171]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9307 (.A([213]), .Y([215]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9308 (.A([44]), .Y([456]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9309 (.A([3]), .Y([1002]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9310 (.A([2148]), .Y([1247]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9311 (.A([1368]), .B([2149]), .X([488]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9312 (.A([488]), .Y([690]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9313 (.A([1216]), .B([2150]), .X([2151]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9314 (.A([1316]), .B([1346]), .X([608]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9315 (.A([2151]), .B([608]), .X([666]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9316 (.A([488]), .B([666]), .X([2039]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9317 (.A([1316]), .B([2152]), .X([2153]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9318 (.A([2151]), .B([2153]), .X([2154]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9319 (.A([1383]), .B([2155]), .X([614]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9320 (.A([614]), .Y([1123]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9321 (.A([2154]), .B([614]), .X([1274]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9322 (.A([1274]), .Y([2156]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9323 (.A([2039]), .B([1274]), .Y([1599]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9324 (.A([1368]), .B([1383]), .X([605]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9325 (.A([605]), .Y([2157]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9326 (.A([1216]), .B([1288]), .X([641]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9327 (.A([2153]), .B([641]), .X([1153]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9328 (.A([605]), .B([1153]), .X([1160]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9329 (.A([488]), .B([2154]), .X([1161]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9330 (.A([1288]), .B([2158]), .X([609]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9331 (.A([1346]), .B([2159]), .X([642]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9332 (.A([609]), .B([642]), .X([654]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9333 (.A([488]), .B([654]), .X([1132]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9334 (.A([1161]), .B([1132]), .Y([1264]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9335 (.A([2039]), .B([1160]), .Y([1563]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9336 (.A([2156]), .B([1264]), .X([2160]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9337 (.A([1563]), .B([2160]), .X([603]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9338 (.A([603]), .Y([719]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9339 (.A([2158]), .B([2150]), .X([2161]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9340 (.A([2153]), .B([2161]), .X([623]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9341 (.A([605]), .B([623]), .X([1125]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9342 (.A([2159]), .B([2152]), .X([2162]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9343 (.A([641]), .B([2162]), .X([2163]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9344 (.A([488]), .B([2163]), .X([629]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9345 (.A([1125]), .B([629]), .Y([2164]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9346 (.A([2161]), .B([2162]), .X([606]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9347 (.A([614]), .B([606]), .X([2165]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9348 (.A([2165]), .Y([697]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9349 (.A([488]), .B([1153]), .X([1188]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9350 (.A([2165]), .B([1188]), .Y([634]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9351 (.A([2151]), .B([2162]), .X([489]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9352 (.A([614]), .B([489]), .X([694]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9353 (.A([694]), .Y([1265]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9354 (.A([614]), .B([2163]), .X([1302]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9355 (.A([694]), .B([1302]), .Y([2166]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9356 (.A([2164]), .B([2166]), .X([2167]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9357 (.A([634]), .B([2167]), .X([2168]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9358 (.A([603]), .B([2168]), .X([2169]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9359 (.A([605]), .B([2163]), .X([1066]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9360 (.A([1066]), .Y([472]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9361 (.A([2169]), .B([472]), .X([2170]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9362 (.A([608]), .B([641]), .X([615]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9363 (.A([2155]), .B([2149]), .X([611]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9364 (.A([615]), .B([611]), .X([1133]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9365 (.A([608]), .B([2161]), .X([639]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9366 (.A([614]), .B([639]), .X([617]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9367 (.A([1133]), .B([617]), .Y([1359]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9368 (.A([605]), .B([489]), .X([1130]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9369 (.A([666]), .B([605]), .X([2171]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9370 (.A([1130]), .B([2171]), .Y([1276]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9371 (.A([1359]), .B([1276]), .X([1565]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9372 (.A([1565]), .Y([2172]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9373 (.A([1449]), .B([2172]), .Y([2173]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9374 (.A([2170]), .B([2173]), .X([2174]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9375 (.A([2175]), .B([1565]), .Y([2176]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9376 (.A([1410]), .B([472]), .Y([2177]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9377 (.A([2176]), .B([2177]), .Y([2178]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9378 (.A([2169]), .B([2178]), .X([2179]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9379 (.A([2179]), .Y([2180]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9380 (.A([2174]), .B([2180]), .Y([588]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9381 (.A([588]), .Y([737]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9382 (.A([1274]), .B([1302]), .Y([1335]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9383 (.A([1335]), .Y([1200]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9384 (.A([634]), .B([1335]), .X([1143]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9385 (.A([481]), .B([2181]), .Y([2182]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9386 (.A([1066]), .B([2182]), .X([2183]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9387 (.A([44]), .B([1066]), .Y([2184]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9388 (.A([2183]), .B([2184]), .Y([2185]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9389 (.A([1143]), .B([2185]), .X([2186]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9390 (.A([2164]), .B([2186]), .X([2187]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9391 (.A([39]), .B([2187]), .Y([2188]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9392 (.A([2188]), .Y([2189]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9393 (.A([1422]), .B([2170]), .X([2190]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9394 (.A([1386]), .B([472]), .Y([2191]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9395 (.A([2172]), .B([2191]), .Y([2192]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9396 (.A([2192]), .Y([2193]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9397 (.A([2190]), .B([2193]), .Y([600]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9398 (.A([600]), .Y([593]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9399 (.A([2189]), .B([600]), .Y([2194]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9400 (.A([737]), .B([2194]), .X([2195]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9401 (.A([2196]), .B([2197]), .X([2198]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9402 (.A([2199]), .B([2198]), .X([2200]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9403 (.A([1886]), .B([2196]), .X([2201]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9404 (.A([1923]), .B([2201]), .X([2202]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9405 (.A([2200]), .B([2202]), .Y([2203]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9406 (.A([1923]), .B([2197]), .X([2204]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9407 (.A([1886]), .B([2199]), .X([2205]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9408 (.A([2204]), .B([2205]), .Y([2206]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9409 (.A([2203]), .B([2206]), .X([2207]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9410 (.A([2196]), .B([2207]), .X([2208]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9411 (.A([44]), .B([2208]), .Y([2209]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9412 (.A([263]), .B([2209]), .Y([2210]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9413 (.A([263]), .B([2209]), .X([2211]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9414 (.A([2210]), .B([2211]), .Y([2212]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9415 (.A([1274]), .B([2212]), .Y([2213]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9416 (.A([39]), .B([2214]), .X([2215]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9417 (.A([433]), .B([20]), .X([2216]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9418 (.A([2215]), .B([2216]), .Y([567]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9419 (.A([567]), .Y([256]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9420 (.A([1274]), .B([256]), .X([2217]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9421 (.A([2217]), .Y([2218]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9422 (.A([2189]), .B([2213]), .Y([2219]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9423 (.A([2218]), .B([2219]), .X([2220]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9424 (.A([2195]), .B([2220]), .X([2221]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9425 (.A([597]), .B([2195]), .Y([2222]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9426 (.A([2221]), .B([2222]), .Y([2223]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9427 (.A([286]), .B([2203]), .Y([2224]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9428 (.A([286]), .B([2203]), .X([2225]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9429 (.A([2224]), .B([2225]), .Y([2226]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9430 (.A([2211]), .B([2226]), .Y([2227]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9431 (.A([2211]), .B([2226]), .X([2228]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9432 (.A([2227]), .B([2228]), .Y([2229]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9433 (.A([1274]), .B([2229]), .Y([2230]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9434 (.A([39]), .B([2231]), .X([2232]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9435 (.A([433]), .B([21]), .X([2233]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9436 (.A([2232]), .B([2233]), .Y([508]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9437 (.A([508]), .Y([281]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9438 (.A([1274]), .B([281]), .X([2234]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9439 (.A([2234]), .Y([2235]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9440 (.A([2189]), .B([2230]), .Y([2236]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9441 (.A([2235]), .B([2236]), .X([2237]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9442 (.A([2195]), .B([2237]), .X([2238]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9443 (.A([2134]), .B([2195]), .Y([2239]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9444 (.A([2238]), .B([2239]), .Y([2240]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9445 (.A([2224]), .B([2228]), .Y([2241]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9446 (.A([2241]), .Y([2242]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9447 (.A([309]), .B([2200]), .X([2243]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9448 (.A([309]), .B([2200]), .Y([2244]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9449 (.A([2243]), .B([2244]), .Y([2245]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9450 (.A([2242]), .B([2245]), .Y([2246]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9451 (.A([2242]), .B([2245]), .X([2247]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9452 (.A([2246]), .B([2247]), .Y([2248]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9453 (.A([1274]), .B([2248]), .Y([2249]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9454 (.A([39]), .B([2250]), .X([2251]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9455 (.A([433]), .B([22]), .X([2252]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9456 (.A([2251]), .B([2252]), .Y([1015]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9457 (.A([1015]), .Y([305]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9458 (.A([1274]), .B([305]), .X([2253]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9459 (.A([2189]), .B([2253]), .Y([2254]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9460 (.A([2254]), .Y([2255]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9461 (.A([2249]), .B([2255]), .Y([2256]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9462 (.A([2195]), .B([2256]), .X([2257]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9463 (.A([739]), .B([2195]), .Y([2258]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9464 (.A([2257]), .B([2258]), .Y([2259]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9465 (.A([2243]), .B([2247]), .Y([2260]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9466 (.A([145]), .B([2202]), .Y([2261]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9467 (.A([145]), .B([2202]), .X([2262]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9468 (.A([2261]), .B([2262]), .Y([2263]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9469 (.A([2263]), .Y([2264]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9470 (.A([2260]), .B([2264]), .Y([2265]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9471 (.A([2260]), .B([2264]), .X([2266]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9472 (.A([2265]), .B([2266]), .Y([2267]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9473 (.A([2156]), .B([2267]), .X([2268]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9474 (.A([39]), .B([2269]), .X([2270]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9475 (.A([433]), .B([23]), .X([2271]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9476 (.A([2270]), .B([2271]), .Y([468]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9477 (.A([468]), .Y([329]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9478 (.A([1274]), .B([329]), .X([2272]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9479 (.A([2189]), .B([2272]), .Y([2273]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9480 (.A([2273]), .Y([2274]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9481 (.A([2268]), .B([2274]), .Y([2275]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9482 (.A([2195]), .B([2275]), .X([2276]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9483 (.A([768]), .B([2195]), .Y([2277]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9484 (.A([2276]), .B([2277]), .Y([2278]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9485 (.A([2279]), .B([2198]), .X([2280]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9486 (.A([550]), .B([2201]), .X([2281]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9487 (.A([2280]), .B([2281]), .Y([2282]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9488 (.A([550]), .B([2197]), .X([2283]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9489 (.A([1886]), .B([2279]), .X([2284]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9490 (.A([2283]), .B([2284]), .Y([2285]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9491 (.A([2282]), .B([2285]), .X([2286]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9492 (.A([2196]), .B([2286]), .X([2287]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9493 (.A([44]), .B([2287]), .Y([2288]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9494 (.A([171]), .B([2288]), .Y([2289]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9495 (.A([171]), .B([2288]), .X([2290]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9496 (.A([2289]), .B([2290]), .Y([2291]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9497 (.A([1274]), .B([2291]), .Y([2292]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9498 (.A([39]), .B([24]), .Y([2293]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9499 (.A([433]), .B([2294]), .Y([2295]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9500 (.A([2293]), .B([2295]), .Y([352]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9501 (.A([1274]), .B([352]), .X([2296]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9502 (.A([2296]), .Y([2297]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9503 (.A([2189]), .B([2292]), .Y([2298]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9504 (.A([2297]), .B([2298]), .X([2299]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9505 (.A([2195]), .B([2299]), .X([2300]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9506 (.A([797]), .B([2195]), .Y([2301]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9507 (.A([2300]), .B([2301]), .Y([2302]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9508 (.A([191]), .B([2282]), .Y([2303]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9509 (.A([191]), .B([2282]), .X([2304]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9510 (.A([2303]), .B([2304]), .Y([2305]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9511 (.A([2290]), .B([2305]), .Y([2306]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9512 (.A([2290]), .B([2305]), .X([2307]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9513 (.A([2306]), .B([2307]), .Y([2308]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9514 (.A([1274]), .B([2308]), .Y([2309]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9515 (.A([39]), .B([2310]), .X([2311]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9516 (.A([433]), .B([25]), .X([2312]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9517 (.A([2311]), .B([2312]), .Y([1028]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9518 (.A([1028]), .Y([375]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9519 (.A([1274]), .B([375]), .X([2313]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9520 (.A([2313]), .Y([2314]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9521 (.A([2189]), .B([2309]), .Y([2315]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9522 (.A([2314]), .B([2315]), .X([2316]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9523 (.A([2195]), .B([2316]), .X([2317]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9524 (.A([826]), .B([2195]), .Y([2318]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9525 (.A([2317]), .B([2318]), .Y([2319]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9526 (.A([2303]), .B([2307]), .Y([2320]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9527 (.A([2320]), .Y([2321]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9528 (.A([215]), .B([2280]), .X([2322]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9529 (.A([215]), .B([2280]), .Y([2323]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9530 (.A([2322]), .B([2323]), .Y([2324]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9531 (.A([2321]), .B([2324]), .Y([2325]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9532 (.A([2321]), .B([2324]), .X([2326]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9533 (.A([2325]), .B([2326]), .Y([2327]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9534 (.A([1274]), .B([2327]), .Y([2328]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9535 (.A([39]), .B([2329]), .X([2330]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9536 (.A([433]), .B([26]), .X([2331]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9537 (.A([2330]), .B([2331]), .Y([1033]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9538 (.A([1033]), .Y([398]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9539 (.A([1274]), .B([398]), .X([2332]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9540 (.A([2189]), .B([2332]), .Y([2333]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9541 (.A([2333]), .Y([2334]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9542 (.A([2328]), .B([2334]), .Y([2335]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9543 (.A([2195]), .B([2335]), .X([2336]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9544 (.A([855]), .B([2195]), .Y([2337]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9545 (.A([2336]), .B([2337]), .Y([2338]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9546 (.A([2322]), .B([2326]), .Y([2339]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9547 (.A([234]), .B([2281]), .Y([2340]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9548 (.A([234]), .B([2281]), .X([2341]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9549 (.A([2340]), .B([2341]), .Y([2342]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9550 (.A([2339]), .B([2342]), .X([2343]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9551 (.A([2339]), .B([2342]), .Y([2344]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9552 (.A([2343]), .B([2344]), .Y([2345]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9553 (.A([1274]), .B([2345]), .Y([2346]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9554 (.A([433]), .B([2347]), .Y([2348]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9555 (.A([39]), .B([27]), .Y([585]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9556 (.A([2348]), .B([585]), .Y([419]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9557 (.A([1274]), .B([419]), .X([2349]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9558 (.A([2189]), .B([2349]), .Y([2350]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9559 (.A([2350]), .Y([2351]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9560 (.A([2346]), .B([2351]), .Y([2352]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9561 (.A([2195]), .B([2352]), .X([2353]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9562 (.A([884]), .B([2195]), .Y([2354]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9563 (.A([2353]), .B([2354]), .Y([2355]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9564 (.A([588]), .B([2194]), .X([2356]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9565 (.A([2135]), .B([2356]), .Y([2357]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9566 (.A([2220]), .B([2356]), .X([2358]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9567 (.A([2357]), .B([2358]), .Y([2359]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9568 (.A([707]), .B([2356]), .Y([2360]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9569 (.A([2237]), .B([2356]), .X([2361]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9570 (.A([2360]), .B([2361]), .Y([2362]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9571 (.A([736]), .B([2356]), .Y([2363]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9572 (.A([2256]), .B([2356]), .X([2364]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9573 (.A([2363]), .B([2364]), .Y([2365]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9574 (.A([2275]), .B([2356]), .X([2366]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9575 (.A([766]), .B([2356]), .Y([2367]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9576 (.A([2366]), .B([2367]), .Y([2368]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9577 (.A([2299]), .B([2356]), .X([2369]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9578 (.A([795]), .B([2356]), .Y([2370]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9579 (.A([2369]), .B([2370]), .Y([2371]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9580 (.A([2316]), .B([2356]), .X([2372]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9581 (.A([824]), .B([2356]), .Y([2373]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9582 (.A([2372]), .B([2373]), .Y([2374]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9583 (.A([2335]), .B([2356]), .X([2375]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9584 (.A([853]), .B([2356]), .Y([2376]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9585 (.A([2375]), .B([2376]), .Y([2377]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9586 (.A([882]), .B([2356]), .Y([2378]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9587 (.A([2352]), .B([2356]), .X([2379]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9588 (.A([2378]), .B([2379]), .Y([2380]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9589 (.A([588]), .B([593]), .Y([482]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9590 (.A([2188]), .B([482]), .X([2381]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9591 (.A([590]), .B([2381]), .Y([2382]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9592 (.A([2220]), .B([2381]), .X([2383]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9593 (.A([2382]), .B([2383]), .Y([2384]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9594 (.A([2237]), .B([2381]), .X([2385]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9595 (.A([711]), .B([2381]), .Y([2386]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9596 (.A([2385]), .B([2386]), .Y([2387]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9597 (.A([743]), .B([2381]), .Y([2388]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9598 (.A([2256]), .B([2381]), .X([2389]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9599 (.A([2388]), .B([2389]), .Y([2390]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9600 (.A([2275]), .B([2381]), .X([2391]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9601 (.A([775]), .B([2381]), .Y([2392]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9602 (.A([2391]), .B([2392]), .Y([2393]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9603 (.A([801]), .B([2381]), .Y([2394]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9604 (.A([2299]), .B([2381]), .X([2395]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9605 (.A([2394]), .B([2395]), .Y([2396]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9606 (.A([2316]), .B([2381]), .X([2397]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9607 (.A([830]), .B([2381]), .Y([2398]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9608 (.A([2397]), .B([2398]), .Y([2399]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9609 (.A([2335]), .B([2381]), .X([2400]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9610 (.A([859]), .B([2381]), .Y([2401]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9611 (.A([2400]), .B([2401]), .Y([2402]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9612 (.A([2352]), .B([2381]), .X([2403]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9613 (.A([891]), .B([2381]), .Y([2404]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9614 (.A([2403]), .B([2404]), .Y([2405]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9615 (.A([588]), .B([600]), .X([715]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9616 (.A([2188]), .B([715]), .X([2406]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9617 (.A([2136]), .B([2406]), .Y([2407]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9618 (.A([2220]), .B([2406]), .X([2408]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9619 (.A([2407]), .B([2408]), .Y([2409]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9620 (.A([2237]), .B([2406]), .X([2410]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9621 (.A([714]), .B([2406]), .Y([2411]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9622 (.A([2410]), .B([2411]), .Y([2412]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9623 (.A([2256]), .B([2406]), .X([2413]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9624 (.A([746]), .B([2406]), .Y([2414]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9625 (.A([2413]), .B([2414]), .Y([2415]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9626 (.A([772]), .B([2406]), .Y([2416]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9627 (.A([2275]), .B([2406]), .X([2417]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9628 (.A([2416]), .B([2417]), .Y([2418]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9629 (.A([2299]), .B([2406]), .X([2419]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9630 (.A([804]), .B([2406]), .Y([2420]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9631 (.A([2419]), .B([2420]), .Y([2421]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9632 (.A([2316]), .B([2406]), .X([2422]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9633 (.A([833]), .B([2406]), .Y([2423]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9634 (.A([2422]), .B([2423]), .Y([2424]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9635 (.A([2335]), .B([2406]), .X([2425]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9636 (.A([862]), .B([2406]), .Y([2426]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9637 (.A([2425]), .B([2426]), .Y([2427]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9638 (.A([888]), .B([2406]), .Y([2428]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9639 (.A([2352]), .B([2406]), .X([2429]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9640 (.A([2428]), .B([2429]), .Y([2430]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9641 (.A([1963]), .B([550]), .X([2431]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9642 (.A([1963]), .B([550]), .Y([2432]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9643 (.A([2431]), .B([2432]), .Y([2433]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9644 (.A([1513]), .B([234]), .Y([2434]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9645 (.A([1513]), .B([234]), .X([2435]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9646 (.A([2434]), .B([2435]), .Y([2436]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9647 (.A([2433]), .B([2436]), .Y([2437]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9648 (.A([2433]), .B([2436]), .X([2438]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9649 (.A([2437]), .B([2438]), .Y([2439]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9650 (.A([2139]), .B([546]), .Y([2440]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9651 (.A([2440]), .Y([2441]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9652 (.A([2439]), .B([2441]), .Y([2442]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9653 (.A([2138]), .B([456]), .Y([2443]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9654 (.A([2137]), .B([2443]), .Y([2444]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9655 (.A([2444]), .Y([2445]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9656 (.A([2442]), .B([2445]), .Y([2446]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9657 (.A([2446]), .Y([2447]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9658 (.A([462]), .B([213]), .Y([2448]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9659 (.A([642]), .B([2161]), .X([2449]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9660 (.A([488]), .B([2449]), .X([469]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9661 (.A([469]), .Y([542]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9662 (.A([472]), .B([469]), .Y([2450]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9663 (.A([2450]), .Y([466]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9664 (.A([2448]), .B([466]), .Y([2451]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9665 (.A([2447]), .B([2451]), .X([2452]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9666 (.A([609]), .B([2162]), .X([2453]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9667 (.A([605]), .B([2453]), .X([1113]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9668 (.A([1113]), .Y([1517]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9669 (.A([511]), .B([1517]), .Y([2454]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9670 (.A([472]), .B([2454]), .X([494]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9671 (.A([469]), .B([494]), .Y([2455]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9672 (.A([2455]), .Y([501]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9673 (.A([2137]), .B([1066]), .X([476]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9674 (.A([2138]), .B([546]), .X([2456]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9675 (.A([462]), .B([2456]), .X([2457]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9676 (.A([472]), .B([2457]), .Y([2458]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9677 (.A([1254]), .B([2458]), .Y([2459]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9678 (.A([501]), .B([2459]), .Y([2460]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9679 (.A([398]), .B([2455]), .Y([2461]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9680 (.A([2460]), .B([2461]), .Y([2462]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9681 (.A([2452]), .B([2462]), .Y([2463]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9682 (.A([2463]), .Y([2464]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9683 (.A([433]), .B([1066]), .X([1404]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9684 (.A([1404]), .Y([1387]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9685 (.A([462]), .B([1404]), .Y([2465]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9686 (.A([2000]), .B([398]), .X([2466]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9687 (.A([37]), .B([2467]), .Y([2468]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9688 (.A([1988]), .B([37]), .X([2092]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9689 (.A([1988]), .B([2467]), .X([2469]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9690 (.A([2092]), .B([2469]), .Y([2470]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9691 (.A([1983]), .B([2468]), .Y([2471]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9692 (.A([2000]), .B([2145]), .Y([2472]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9693 (.A([2466]), .B([2472]), .Y([2473]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9694 (.A([2471]), .B([2473]), .X([2474]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9695 (.A([2474]), .Y([2475]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9696 (.A([2000]), .B([419]), .X([2476]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9697 (.A([2000]), .B([2146]), .Y([2477]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9698 (.A([2470]), .B([2477]), .Y([2478]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9699 (.A([2478]), .Y([2479]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9700 (.A([2476]), .B([2479]), .Y([1455]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9701 (.A([1455]), .Y([2480]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9702 (.A([2000]), .B([352]), .X([2481]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9703 (.A([2000]), .B([2144]), .Y([2482]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9704 (.A([2481]), .B([2482]), .Y([2483]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9705 (.A([2471]), .B([2483]), .X([1349]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9706 (.A([1349]), .Y([1174]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9707 (.A([44]), .B([2471]), .Y([2484]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9708 (.A([1349]), .B([2484]), .Y([1094]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9709 (.A([1094]), .Y([1058]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9710 (.A([1455]), .B([2484]), .Y([450]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9711 (.A([450]), .Y([1497]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9712 (.A([1349]), .B([1497]), .Y([1087]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9713 (.A([1087]), .Y([1083]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9714 (.A([2000]), .B([1028]), .X([2485]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9715 (.A([2000]), .B([1026]), .Y([2486]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9716 (.A([2485]), .B([2486]), .Y([2487]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9717 (.A([2470]), .B([2487]), .Y([1506]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9718 (.A([1094]), .B([1506]), .X([1049]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9719 (.A([1087]), .B([1506]), .X([1046]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9720 (.A([2474]), .B([2484]), .Y([445]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9721 (.A([1046]), .B([445]), .X([1040]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9722 (.A([2000]), .B([281]), .X([2488]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9723 (.A([2000]), .B([2141]), .Y([2489]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9724 (.A([2470]), .B([2489]), .Y([2490]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9725 (.A([2490]), .Y([2491]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9726 (.A([2488]), .B([2491]), .Y([2492]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9727 (.A([2492]), .Y([2493]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9728 (.A([2000]), .B([256]), .X([2494]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9729 (.A([2000]), .B([2140]), .Y([2495]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9730 (.A([2494]), .B([2495]), .Y([2496]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9731 (.A([2471]), .B([2496]), .X([2497]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9732 (.A([2497]), .Y([1097]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9733 (.A([2484]), .B([2497]), .Y([2498]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9734 (.A([2493]), .B([2498]), .X([1055]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9735 (.A([1055]), .Y([1431]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9736 (.A([2000]), .B([329]), .X([2499]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9737 (.A([2000]), .B([2143]), .Y([2500]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9738 (.A([2499]), .B([2500]), .Y([2501]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9739 (.A([2471]), .B([2501]), .X([2502]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9740 (.A([2000]), .B([305]), .X([2503]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9741 (.A([2000]), .B([2142]), .Y([2504]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9742 (.A([2470]), .B([2504]), .Y([2505]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9743 (.A([2505]), .Y([2506]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9744 (.A([2503]), .B([2506]), .Y([1061]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9745 (.A([2484]), .B([1061]), .Y([1069]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9746 (.A([2502]), .B([1069]), .X([1395]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9747 (.A([1055]), .B([1395]), .X([1047]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9748 (.A([1404]), .B([1047]), .X([2507]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9749 (.A([1040]), .B([2507]), .X([2508]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9750 (.A([2465]), .B([2508]), .Y([2509]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9751 (.A([2043]), .B([1404]), .Y([2510]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9752 (.A([1083]), .B([1506]), .Y([1076]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9753 (.A([2475]), .B([1076]), .X([1101]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9754 (.A([2507]), .B([1101]), .X([2511]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9755 (.A([2510]), .B([2511]), .Y([2512]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9756 (.A([554]), .B([1404]), .Y([2513]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9757 (.A([2474]), .B([1497]), .Y([1460]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9758 (.A([2484]), .B([1506]), .Y([440]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9759 (.A([440]), .Y([2514]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9760 (.A([1349]), .B([440]), .X([1412]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9761 (.A([2507]), .B([1412]), .X([2515]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9762 (.A([1460]), .B([2515]), .X([2516]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9763 (.A([2513]), .B([2516]), .Y([2517]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9764 (.A([552]), .B([1404]), .Y([2518]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9765 (.A([1094]), .B([440]), .Y([2519]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9766 (.A([2507]), .B([2519]), .X([2520]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9767 (.A([1460]), .B([2520]), .X([2521]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9768 (.A([2518]), .B([2521]), .Y([2522]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9769 (.A([453]), .B([1404]), .Y([2523]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9770 (.A([450]), .B([445]), .Y([1477]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9771 (.A([2515]), .B([1477]), .X([2524]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9772 (.A([2523]), .B([2524]), .Y([2525]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9773 (.A([454]), .B([1404]), .Y([2526]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9774 (.A([2520]), .B([1477]), .X([2527]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9775 (.A([2526]), .B([2527]), .Y([2528]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9776 (.A([2021]), .B([1404]), .Y([2529]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9777 (.A([2474]), .B([450]), .X([1050]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9778 (.A([2515]), .B([1050]), .X([2530]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9779 (.A([2529]), .B([2530]), .Y([2531]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9780 (.A([2014]), .B([1404]), .Y([2532]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9781 (.A([2520]), .B([1050]), .X([2533]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9782 (.A([2532]), .B([2533]), .Y([2534]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9783 (.A([2138]), .B([1404]), .Y([2535]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9784 (.A([1455]), .B([445]), .X([1413]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9785 (.A([1413]), .Y([2536]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9786 (.A([2520]), .B([1413]), .X([2537]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9787 (.A([2535]), .B([2537]), .Y([2538]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9788 (.A([511]), .B([1404]), .Y([2539]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9789 (.A([2498]), .B([1061]), .X([2540]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9790 (.A([1055]), .B([1061]), .X([2541]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9791 (.A([1040]), .B([2541]), .X([1463]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9792 (.A([1404]), .B([1463]), .X([2542]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9793 (.A([2539]), .B([2542]), .Y([2543]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9794 (.A([1523]), .B([1404]), .Y([2544]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9795 (.A([2492]), .B([2498]), .X([1072]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9796 (.A([1395]), .B([1072]), .X([1085]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9797 (.A([1061]), .B([1072]), .X([2545]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9798 (.A([1085]), .B([2545]), .Y([2546]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9799 (.A([1404]), .B([450]), .X([2547]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9800 (.A([2547]), .Y([2548]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9801 (.A([2546]), .B([2548]), .Y([2549]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9802 (.A([2514]), .B([2549]), .X([2550]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9803 (.A([450]), .B([1085]), .X([2551]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9804 (.A([2544]), .B([2550]), .Y([2552]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9805 (.A([1050]), .B([1072]), .X([1464]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9806 (.A([1404]), .B([1464]), .X([2553]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9807 (.A([1555]), .B([1404]), .Y([2554]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9808 (.A([2553]), .B([2554]), .Y([2555]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9809 (.A([2484]), .B([2502]), .Y([1062]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9810 (.A([1062]), .Y([2556]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9811 (.A([2541]), .B([2556]), .X([1052]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9812 (.A([1052]), .Y([1043]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9813 (.A([1455]), .B([1094]), .X([1041]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9814 (.A([2474]), .B([1041]), .X([2557]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9815 (.A([1052]), .B([2557]), .X([2558]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9816 (.A([1055]), .B([1477]), .X([1393]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9817 (.A([1174]), .B([1062]), .X([2559]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9818 (.A([1393]), .B([2559]), .X([2560]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9819 (.A([2558]), .B([2560]), .Y([1484]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9820 (.A([2492]), .B([1097]), .Y([1073]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9821 (.A([2475]), .B([1506]), .Y([1088]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9822 (.A([1073]), .B([1088]), .X([1495]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9823 (.A([1497]), .B([1495]), .X([2561]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9824 (.A([1387]), .B([2561]), .Y([2562]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9825 (.A([1484]), .B([2562]), .X([2563]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9826 (.A([484]), .B([1404]), .Y([2564]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9827 (.A([2563]), .B([2564]), .Y([2565]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9828 (.A([2565]), .Y([2566]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9829 (.A([539]), .B([1404]), .Y([2567]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9830 (.A([2549]), .B([2567]), .Y([2568]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9831 (.A([1160]), .B([1066]), .Y([2569]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9832 (.A([39]), .B([2569]), .Y([2570]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9833 (.A([546]), .B([2570]), .Y([2571]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9834 (.A([445]), .B([440]), .Y([1456]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9835 (.A([1073]), .B([2570]), .X([2572]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9836 (.A([1456]), .B([2572]), .X([2573]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9837 (.A([2571]), .B([2573]), .Y([2574]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9838 (.A([1886]), .B([2570]), .Y([2575]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9839 (.A([474]), .B([1497]), .Y([2576]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9840 (.A([2573]), .B([2576]), .X([2577]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9841 (.A([2575]), .B([2577]), .Y([2578]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9842 (.A([1477]), .B([2545]), .X([1473]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9843 (.A([2514]), .B([1473]), .X([2579]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9844 (.A([1047]), .B([2557]), .X([2580]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9845 (.A([2579]), .B([2580]), .Y([2581]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9846 (.A([1387]), .B([2581]), .Y([2582]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9847 (.A([1543]), .B([1404]), .Y([2583]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9848 (.A([2582]), .B([2583]), .Y([2584]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9849 (.A([1506]), .B([1413]), .X([1397]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9850 (.A([1404]), .B([1397]), .X([2585]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9851 (.A([1525]), .B([1404]), .Y([2586]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9852 (.A([2585]), .B([2586]), .Y([2587]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9853 (.A([1196]), .B([1404]), .Y([2588]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9854 (.A([1387]), .B([1413]), .Y([2589]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9855 (.A([2545]), .B([2589]), .X([2590]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9856 (.A([2588]), .B([2590]), .Y([2591]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9857 (.A([2540]), .B([1073]), .Y([2592]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9858 (.A([1193]), .B([1404]), .Y([2593]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9859 (.A([2536]), .B([2592]), .Y([2594]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9860 (.A([1404]), .B([440]), .X([2595]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9861 (.A([2594]), .B([2595]), .X([2596]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9862 (.A([2593]), .B([2596]), .Y([2597]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9863 (.A([1061]), .B([2556]), .Y([1056]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9864 (.A([1073]), .B([1056]), .X([1064]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9865 (.A([1058]), .B([1064]), .X([1219]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9866 (.A([1395]), .B([1073]), .X([1095]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9867 (.A([1387]), .B([1095]), .Y([2598]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9868 (.A([1413]), .B([1072]), .X([2599]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9869 (.A([2599]), .Y([1438]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9870 (.A([1349]), .B([1413]), .X([2600]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9871 (.A([2545]), .B([2600]), .X([2601]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9872 (.A([1219]), .B([2601]), .Y([2602]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9873 (.A([2598]), .B([2602]), .X([2603]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9874 (.A([2175]), .B([1387]), .X([2604]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9875 (.A([2603]), .B([2604]), .Y([2605]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9876 (.A([2605]), .Y([2606]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9877 (.A([481]), .B([1387]), .X([2607]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9878 (.A([1047]), .B([2551]), .Y([2608]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9879 (.A([1058]), .B([2608]), .Y([2609]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9880 (.A([2609]), .Y([2610]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9881 (.A([2540]), .B([1085]), .Y([2611]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9882 (.A([1349]), .B([1397]), .X([1445]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9883 (.A([1097]), .B([1413]), .X([2612]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9884 (.A([2502]), .B([440]), .X([1436]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9885 (.A([1069]), .B([1436]), .X([2613]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9886 (.A([2480]), .B([1506]), .Y([2614]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9887 (.A([2614]), .Y([2615]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9888 (.A([1094]), .B([2614]), .X([1389]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9889 (.A([1041]), .B([1088]), .X([1428]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9890 (.A([1085]), .B([1428]), .X([1479]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9891 (.A([1479]), .Y([1406]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9892 (.A([1073]), .B([2615]), .X([2616]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9893 (.A([1445]), .B([1479]), .Y([2617]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9894 (.A([2611]), .B([2617]), .Y([2618]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9895 (.A([1413]), .B([2613]), .X([2619]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9896 (.A([2498]), .B([2619]), .X([2620]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9897 (.A([2616]), .B([2620]), .Y([2621]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9898 (.A([2621]), .Y([2622]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9899 (.A([2618]), .B([2622]), .Y([2623]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9900 (.A([1049]), .B([2612]), .X([2624]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9901 (.A([1387]), .B([2624]), .Y([2625]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9902 (.A([2623]), .B([2625]), .X([2626]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9903 (.A([2610]), .B([2626]), .X([2627]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9904 (.A([2607]), .B([2627]), .Y([2628]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9905 (.A([2628]), .Y([2629]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9906 (.A([1066]), .B([2471]), .X([2630]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9907 (.A([2151]), .B([642]), .X([621]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9908 (.A([605]), .B([621]), .X([172]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9909 (.A([172]), .Y([148]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9910 (.A([583]), .B([550]), .X([2631]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9911 (.A([583]), .B([550]), .Y([2632]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9912 (.A([2631]), .B([2632]), .Y([1184]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9913 (.A([148]), .B([1184]), .Y([1331]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9914 (.A([2630]), .B([1331]), .Y([2633]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9915 (.A([1125]), .B([1113]), .Y([2634]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9916 (.A([605]), .B([2449]), .X([264]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9917 (.A([264]), .Y([287]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9918 (.A([488]), .B([2453]), .X([2635]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9919 (.A([264]), .B([2635]), .Y([2636]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9920 (.A([2634]), .B([2636]), .X([2637]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9921 (.A([2633]), .B([2637]), .X([2638]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9922 (.A([44]), .B([172]), .Y([1578]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9923 (.A([472]), .B([1578]), .X([2639]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9924 (.A([2639]), .Y([2640]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9925 (.A([614]), .B([2449]), .X([2641]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9926 (.A([2153]), .B([609]), .X([631]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9927 (.A([488]), .B([631]), .X([2642]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9928 (.A([2641]), .B([2642]), .Y([1115]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9929 (.A([614]), .B([631]), .X([1126]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9930 (.A([1126]), .Y([2643]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9931 (.A([1115]), .B([2643]), .X([650]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9932 (.A([605]), .B([654]), .X([1295]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9933 (.A([1295]), .Y([1262]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9934 (.A([666]), .B([615]), .Y([691]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9935 (.A([2157]), .B([691]), .Y([1201]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9936 (.A([1295]), .B([1201]), .Y([1144]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9937 (.A([650]), .B([1144]), .X([2644]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9938 (.A([2640]), .B([2644]), .X([2645]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9939 (.A([2638]), .B([2645]), .X([2646]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9940 (.A([614]), .B([2453]), .X([2647]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9941 (.A([2635]), .B([2647]), .Y([1119]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9942 (.A([650]), .B([1119]), .X([146]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9943 (.A([2154]), .B([605]), .X([150]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9944 (.A([150]), .Y([199]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9945 (.A([1066]), .B([172]), .Y([2648]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9946 (.A([199]), .B([2648]), .X([1141]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9947 (.A([287]), .B([1141]), .X([2649]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9948 (.A([146]), .B([2649]), .X([2650]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9949 (.A([2630]), .B([2650]), .Y([254]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9950 (.A([287]), .B([254]), .X([143]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9951 (.A([675]), .B([143]), .Y([2651]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9952 (.A([516]), .B([146]), .Y([2652]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9953 (.A([1066]), .B([2470]), .X([2653]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9954 (.A([2653]), .Y([153]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9955 (.A([678]), .B([153]), .Y([2654]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9956 (.A([263]), .B([172]), .X([681]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9957 (.A([2654]), .B([681]), .Y([2655]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9958 (.A([2655]), .Y([2656]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9959 (.A([2652]), .B([2656]), .Y([2657]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9960 (.A([2657]), .Y([2658]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9961 (.A([2651]), .B([2658]), .Y([2659]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9962 (.A([2646]), .B([2659]), .Y([2660]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9963 (.A([2660]), .Y([2661]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9964 (.A([2646]), .B([2659]), .X([2662]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9965 (.A([2660]), .B([2662]), .Y([2663]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9966 (.A([39]), .B([2663]), .Y([2664]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9967 (.A([675]), .B([39]), .X([2665]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9968 (.A([2664]), .B([2665]), .Y([2666]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9969 (.A([2666]), .Y([2667]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9970 (.A([721]), .B([143]), .Y([2668]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9971 (.A([286]), .B([146]), .Y([2669]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9972 (.A([724]), .B([153]), .Y([2670]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9973 (.A([286]), .B([148]), .Y([2671]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9974 (.A([2671]), .Y([729]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9975 (.A([2672]), .B([199]), .Y([2673]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9976 (.A([2670]), .B([2673]), .Y([2674]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9977 (.A([2669]), .B([2671]), .Y([2675]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9978 (.A([2674]), .B([2675]), .X([2676]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9979 (.A([2676]), .Y([2677]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9980 (.A([2668]), .B([2677]), .Y([2678]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9981 (.A([2661]), .B([2678]), .Y([2679]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9982 (.A([2679]), .Y([132]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9983 (.A([2661]), .B([2678]), .X([2680]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9984 (.A([2679]), .B([2680]), .Y([2681]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9985 (.A([39]), .B([2681]), .Y([2682]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9986 (.A([39]), .B([721]), .X([2683]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9987 (.A([2682]), .B([2683]), .Y([2684]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9988 (.A([2684]), .Y([2685]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9989 (.A([138]), .B([143]), .Y([130]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9990 (.A([518]), .B([146]), .Y([2686]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9991 (.A([2686]), .Y([127]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9992 (.A([753]), .B([153]), .Y([2687]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9993 (.A([309]), .B([172]), .X([2688]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9994 (.A([2688]), .Y([124]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9995 (.A([1531]), .B([1995]), .Y([2689]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9996 (.A([1995]), .B([2690]), .X([2691]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9997 (.A([2689]), .B([2691]), .Y([2692]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9998 (.A([150]), .B([2692]), .X([2693]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9999 (.A([2687]), .B([2693]), .Y([125]));
  sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:40:hilomap_worker$12031 (.HI([2694]));
  sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:40:hilomap_worker$8815 (.HI([60]));
  sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:48:hilomap_worker$8817 (.LO([44]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11708 (.A([531]), .Y([2695]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11709 (.A([577]), .Y([2696]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11710 (.A([2110]), .Y([2697]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11711 (.A([2121]), .Y([2698]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11712 (.A([44]), .Y([2699]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11713 (.A([60]), .Y([2700]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11714 (.A([60]), .Y([2701]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11715 (.A([44]), .Y([2702]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11716 (.A([60]), .Y([2703]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11717 (.A([44]), .Y([2704]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11718 (.A([60]), .Y([2705]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11719 (.A([60]), .Y([2706]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11720 (.A([44]), .Y([2707]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11721 (.A([60]), .Y([2708]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11722 (.A([44]), .Y([2709]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11723 (.A([44]), .Y([2710]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11724 (.A([44]), .Y([2711]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11725 (.A([60]), .Y([2712]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11726 (.A([44]), .Y([2713]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11727 (.A([60]), .Y([2714]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11728 (.A([44]), .Y([2715]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11729 (.A([44]), .Y([2716]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11730 (.A([60]), .Y([2717]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11731 (.A([44]), .Y([2718]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11732 (.A([44]), .Y([2719]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11733 (.A([60]), .Y([2720]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11734 (.A([44]), .Y([2721]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11735 (.A([44]), .Y([2722]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11736 (.A([60]), .Y([2723]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11737 (.A([44]), .Y([2724]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11738 (.A([44]), .Y([2725]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11739 (.A([60]), .Y([2726]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11740 (.A([60]), .Y([2727]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11741 (.A([44]), .Y([2728]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11742 (.A([44]), .Y([2729]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11743 (.A([44]), .Y([2730]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11744 (.A([60]), .Y([2731]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11745 (.A([60]), .Y([2732]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11746 (.A([44]), .Y([2733]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11747 (.A([44]), .Y([2734]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11748 (.A([60]), .Y([2735]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11749 (.A([60]), .Y([2736]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11750 (.A([60]), .Y([2737]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11751 (.A([44]), .Y([2738]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11752 (.A([60]), .Y([2739]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11753 (.A([44]), .Y([2740]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11754 (.A([2741]), .Y([2742]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11755 (.A([60]), .Y([2743]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11756 (.A([44]), .Y([2744]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11757 (.A([44]), .Y([2745]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11758 (.A([44]), .Y([2746]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11759 (.A([60]), .Y([2747]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11760 (.A([44]), .Y([2748]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11761 (.A([44]), .Y([2749]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11762 (.A([60]), .Y([2750]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11763 (.A([44]), .Y([2751]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11764 (.A([60]), .Y([2752]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11765 (.A([60]), .Y([2753]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11766 (.A([44]), .Y([2754]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11767 (.A([44]), .Y([2755]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11768 (.A([60]), .Y([2756]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11769 (.A([44]), .Y([2757]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11770 (.A([60]), .Y([2758]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11771 (.A([60]), .Y([2759]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11772 (.A([44]), .Y([2760]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11773 (.A([60]), .Y([2761]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11774 (.A([44]), .Y([2762]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11775 (.A([44]), .Y([2763]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11776 (.A([60]), .Y([2764]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11777 (.A([60]), .Y([2765]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11778 (.A([44]), .Y([2766]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11779 (.A([60]), .Y([2767]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11780 (.A([60]), .Y([2768]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11781 (.A([60]), .Y([2769]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11782 (.A([44]), .Y([2770]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11783 (.A([60]), .Y([2771]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11784 (.A([44]), .Y([2772]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11785 (.A([60]), .Y([2773]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11786 (.A([60]), .Y([2774]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11787 (.A([44]), .Y([2775]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11788 (.A([44]), .Y([2776]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11789 (.A([60]), .Y([2777]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11790 (.A([44]), .Y([2778]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11791 (.A([60]), .Y([2779]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11792 (.A([44]), .Y([2780]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11793 (.A([44]), .Y([2781]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11794 (.A([44]), .Y([2782]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11795 (.A([60]), .Y([2783]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11796 (.A([44]), .Y([2784]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11797 (.A([60]), .Y([2785]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11798 (.A([60]), .Y([2786]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11799 (.A([60]), .Y([2787]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11800 (.A([60]), .Y([2788]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11801 (.A([44]), .Y([2789]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11802 (.A([44]), .Y([2790]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11803 (.A([60]), .Y([2791]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11804 (.A([44]), .Y([2792]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11805 (.A([60]), .Y([2793]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11806 (.A([60]), .Y([2794]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11807 (.A([44]), .Y([2795]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11808 (.A([44]), .Y([2796]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11809 (.A([60]), .Y([2797]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11810 (.A([60]), .Y([2798]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11811 (.A([44]), .Y([2799]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11812 (.A([60]), .Y([2800]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11813 (.A([60]), .Y([2801]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11814 (.A([60]), .Y([2802]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11815 (.A([44]), .Y([2803]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11816 (.A([44]), .Y([2804]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11817 (.A([44]), .Y([2805]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11818 (.A([60]), .Y([2806]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11819 (.A([60]), .Y([2807]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11820 (.A([60]), .Y([2808]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11821 (.A([44]), .Y([2809]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11822 (.A([60]), .Y([2810]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11823 (.A([60]), .Y([2811]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11824 (.A([44]), .Y([2812]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11825 (.A([60]), .Y([2813]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11826 (.A([60]), .Y([2814]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11827 (.A([44]), .Y([2815]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11828 (.A([44]), .Y([2816]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11829 (.A([44]), .Y([2817]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11830 (.A([44]), .Y([2818]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11831 (.A([44]), .Y([2819]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11832 (.A([44]), .Y([2820]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11833 (.A([60]), .Y([2821]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11834 (.A([60]), .Y([2822]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11835 (.A([60]), .Y([2823]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11836 (.A([60]), .Y([2824]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11837 (.A([60]), .Y([2825]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11838 (.A([60]), .Y([2826]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11839 (.A([44]), .Y([2827]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11840 (.A([44]), .Y([2828]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11841 (.A([60]), .Y([2829]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11842 (.A([44]), .Y([2830]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11843 (.A([44]), .Y([2831]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11844 (.A([44]), .Y([2832]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11845 (.A([60]), .Y([2833]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11846 (.A([44]), .Y([2834]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11847 (.A([60]), .Y([2835]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11848 (.A([60]), .Y([2836]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11849 (.A([60]), .Y([2837]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11850 (.A([44]), .Y([2838]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11851 (.A([60]), .Y([2839]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11852 (.A([60]), .Y([2840]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11853 (.A([44]), .Y([2841]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11854 (.A([60]), .Y([2842]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11855 (.A([44]), .Y([2843]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11856 (.A([44]), .Y([2844]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11857 (.A([44]), .Y([2845]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11858 (.A([60]), .Y([2846]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11859 (.A([44]), .Y([2847]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11860 (.A([60]), .Y([2848]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11861 (.A([44]), .Y([2849]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11862 (.A([60]), .Y([2850]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11863 (.A([60]), .Y([2851]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11864 (.A([44]), .Y([2852]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11865 (.A([44]), .Y([2853]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11866 (.A([60]), .Y([2854]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11867 (.A([44]), .Y([2855]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11868 (.A([60]), .Y([2856]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11869 (.A([44]), .Y([2857]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11870 (.A([44]), .Y([2858]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11871 (.A([44]), .Y([2859]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11872 (.A([60]), .Y([2860]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11873 (.A([44]), .Y([2861]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11874 (.A([44]), .Y([2862]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11875 (.A([44]), .Y([2863]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11876 (.A([44]), .Y([2864]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11877 (.A([44]), .Y([2865]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11878 (.A([60]), .Y([2866]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11879 (.A([44]), .Y([2867]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11880 (.A([60]), .Y([2868]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11881 (.A([60]), .Y([2869]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11882 (.A([60]), .Y([2870]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11883 (.A([60]), .Y([2871]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11884 (.A([44]), .Y([2872]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11885 (.A([44]), .Y([2873]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11886 (.A([60]), .Y([2874]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11887 (.A([1196]), .Y([2875]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11888 (.A([562]), .Y([2876]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11889 (.A([44]), .Y([2877]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11890 (.A([1196]), .Y([2878]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11891 (.A([2879]), .Y([2880]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11892 (.A([44]), .Y([2881]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11893 (.A([60]), .Y([2882]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11894 (.A([44]), .Y([2883]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11895 (.A([44]), .Y([2884]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11896 (.A([60]), .Y([2885]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11897 (.A([60]), .Y([2886]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11898 (.A([44]), .Y([2887]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11899 (.A([44]), .Y([2888]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11900 (.A([44]), .Y([2889]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11901 (.A([44]), .Y([2890]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11902 (.A([60]), .Y([2891]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11903 (.A([44]), .Y([2892]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11904 (.A([44]), .Y([2893]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11905 (.A([44]), .Y([2894]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11906 (.A([44]), .Y([2895]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11907 (.A([44]), .Y([2896]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11908 (.A([60]), .Y([2897]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11909 (.A([44]), .Y([2898]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11910 (.A([44]), .Y([2899]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11911 (.A([44]), .Y([2900]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11912 (.A([60]), .Y([2901]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11913 (.A([60]), .Y([2902]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11914 (.A([44]), .Y([2903]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11915 (.A([60]), .Y([2904]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11916 (.A([60]), .Y([2905]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11917 (.A([60]), .Y([2906]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11918 (.A([60]), .Y([2907]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11919 (.A([60]), .Y([2908]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11920 (.A([60]), .Y([2909]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11921 (.A([60]), .Y([2910]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11922 (.A([60]), .Y([2911]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11923 (.A([60]), .Y([2912]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11924 (.A([60]), .Y([2913]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11925 (.A([60]), .Y([2914]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11926 (.A([60]), .Y([2915]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11927 (.A([60]), .Y([2916]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11928 (.A([675]), .Y([2917]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11929 (.A([721]), .Y([2918]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11930 (.A([138]), .Y([2919]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11931 (.A([142]), .Y([2920]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11932 (.A([167]), .Y([2921]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11933 (.A([189]), .Y([2922]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11934 (.A([211]), .Y([2923]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11935 (.A([232]), .Y([2924]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11936 (.A([516]), .Y([2925]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11937 (.A([286]), .Y([2926]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11938 (.A([518]), .Y([2927]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11939 (.A([145]), .Y([2928]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11940 (.A([169]), .Y([2929]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11941 (.A([191]), .Y([2930]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11942 (.A([213]), .Y([2931]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11943 (.A([234]), .Y([2932]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11944 (.A([516]), .Y([2933]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11945 (.A([286]), .Y([2934]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11946 (.A([518]), .Y([2935]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11947 (.A([145]), .Y([2936]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11948 (.A([169]), .Y([2937]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11949 (.A([191]), .Y([2938]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11950 (.A([213]), .Y([2939]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11951 (.A([234]), .Y([2940]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11952 (.A([258]), .Y([2941]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11953 (.A([283]), .Y([2942]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11954 (.A([307]), .Y([2943]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11955 (.A([331]), .Y([2944]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11956 (.A([355]), .Y([2945]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11957 (.A([378]), .Y([2946]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11958 (.A([400]), .Y([2947]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11959 (.A([421]), .Y([2948]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11960 (.A([516]), .Y([2949]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11961 (.A([286]), .Y([2950]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11962 (.A([518]), .Y([2951]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11963 (.A([145]), .Y([2952]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11964 (.A([169]), .Y([2953]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11965 (.A([191]), .Y([2954]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11966 (.A([213]), .Y([2955]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11967 (.A([234]), .Y([2956]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11968 (.A([256]), .Y([2957]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11969 (.A([281]), .Y([2958]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11970 (.A([305]), .Y([2959]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11971 (.A([329]), .Y([2960]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11972 (.A([352]), .Y([2961]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11973 (.A([375]), .Y([2962]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11974 (.A([398]), .Y([2963]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11975 (.A([419]), .Y([2964]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11976 (.A([234]), .Y([2965]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11977 (.A([44]), .Y([45]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11978 (.A([44]), .Y([54]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11979 (.A([44]), .Y([55]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11980 (.A([44]), .Y([56]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11981 (.A([44]), .Y([57]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11982 (.A([44]), .Y([58]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11983 (.A([44]), .Y([59]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11984 (.A([60]), .Y([61]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11985 (.A([60]), .Y([62]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11986 (.A([60]), .Y([63]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11987 (.A([44]), .Y([46]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11988 (.A([60]), .Y([64]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11989 (.A([60]), .Y([65]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11990 (.A([60]), .Y([66]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11991 (.A([60]), .Y([67]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11992 (.A([44]), .Y([68]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11993 (.A([44]), .Y([69]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11994 (.A([44]), .Y([70]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11995 (.A([44]), .Y([71]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11996 (.A([44]), .Y([72]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11997 (.A([44]), .Y([73]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11998 (.A([44]), .Y([47]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11999 (.A([44]), .Y([74]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12000 (.A([44]), .Y([75]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12001 (.A([44]), .Y([76]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12002 (.A([60]), .Y([77]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12003 (.A([60]), .Y([78]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12004 (.A([60]), .Y([79]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12005 (.A([60]), .Y([80]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12006 (.A([60]), .Y([81]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12007 (.A([60]), .Y([82]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12008 (.A([60]), .Y([83]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12009 (.A([44]), .Y([48]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12010 (.A([44]), .Y([49]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12011 (.A([44]), .Y([50]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12012 (.A([44]), .Y([51]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12013 (.A([44]), .Y([52]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12014 (.A([44]), .Y([53]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12015 (.A([44]), .Y([100]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12016 (.A([44]), .Y([101]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12017 (.A([44]), .Y([102]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12018 (.A([44]), .Y([103]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12019 (.A([44]), .Y([104]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12020 (.A([44]), .Y([105]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12021 (.A([44]), .Y([106]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12022 (.A([44]), .Y([107]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12023 (.A([44]), .Y([117]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12024 (.A([44]), .Y([118]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12025 (.A([44]), .Y([119]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12026 (.A([44]), .Y([120]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12027 (.A([44]), .Y([121]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12028 (.A([44]), .Y([122]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12029 (.A([44]), .Y([123]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4105 (.CLK(clk_L0_B0), .D([2223]), .Q([597]), .Q_N([2966]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4106 (.CLK(clk_L0_B0), .D([2240]), .Q([2134]), .Q_N([2967]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4107 (.CLK(clk_L0_B0), .D([2259]), .Q([739]), .Q_N([2968]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4108 (.CLK(clk_L0_B0), .D([2278]), .Q([768]), .Q_N([2969]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4109 (.CLK(clk_L0_B0), .D([2302]), .Q([797]), .Q_N([2970]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4110 (.CLK(clk_L0_B0), .D([2319]), .Q([826]), .Q_N([2971]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4111 (.CLK(clk_L0_B0), .D([2338]), .Q([855]), .Q_N([2972]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4112 (.CLK(clk_L0_B0), .D([2355]), .Q([884]), .Q_N([2973]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4907 (.CLK(clk_L0_B0), .D([2359]), .Q([2135]), .Q_N([2974]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4908 (.CLK(clk_L0_B0), .D([2362]), .Q([707]), .Q_N([2975]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4909 (.CLK(clk_L0_B0), .D([2365]), .Q([736]), .Q_N([2976]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4910 (.CLK(clk_L0_B0), .D([2368]), .Q([766]), .Q_N([2977]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4911 (.CLK(clk_L0_B0), .D([2371]), .Q([795]), .Q_N([2978]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4912 (.CLK(clk_L0_B0), .D([2374]), .Q([824]), .Q_N([2979]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4913 (.CLK(clk_L0_B0), .D([2377]), .Q([853]), .Q_N([2980]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4914 (.CLK(clk_L0_B0), .D([2380]), .Q([882]), .Q_N([2981]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4931 (.CLK(clk_L0_B1), .D([2384]), .Q([590]), .Q_N([2982]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4932 (.CLK(clk_L0_B1), .D([2387]), .Q([711]), .Q_N([2983]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4933 (.CLK(clk_L0_B1), .D([2390]), .Q([743]), .Q_N([2984]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4934 (.CLK(clk_L0_B1), .D([2393]), .Q([775]), .Q_N([2985]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4935 (.CLK(clk_L0_B1), .D([2396]), .Q([801]), .Q_N([2986]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4936 (.CLK(clk_L0_B1), .D([2399]), .Q([830]), .Q_N([2987]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4937 (.CLK(clk_L0_B1), .D([2402]), .Q([859]), .Q_N([2988]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4938 (.CLK(clk_L0_B1), .D([2405]), .Q([891]), .Q_N([2989]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4979 (.CLK(clk_L0_B1), .D([2409]), .Q([2136]), .Q_N([2990]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4980 (.CLK(clk_L0_B1), .D([2412]), .Q([714]), .Q_N([2991]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4981 (.CLK(clk_L0_B1), .D([2415]), .Q([746]), .Q_N([2992]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4982 (.CLK(clk_L0_B1), .D([2418]), .Q([772]), .Q_N([2993]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4983 (.CLK(clk_L0_B1), .D([2421]), .Q([804]), .Q_N([2994]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4984 (.CLK(clk_L0_B1), .D([2424]), .Q([833]), .Q_N([2995]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4985 (.CLK(clk_L0_B1), .D([2427]), .Q([862]), .Q_N([2996]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4986 (.CLK(clk_L0_B1), .D([2430]), .Q([888]), .Q_N([2997]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5134 (.CLK(clk_L0_B2), .D([2464]), .Q([2110]), .Q_N([1251]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5135 (.CLK(clk_L0_B2), .D([1992]), .Q([1988]), .Q_N([2690]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5136 (.CLK(clk_L0_B3), .D([38]), .Q([2998]), .Q_N([1985]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5137 (.CLK(clk_L0_B2), .D([2509]), .Q([462]), .Q_N([2181]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5138 (.CLK(clk_L0_B2), .D([2512]), .Q([2043]), .Q_N([2999]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5139 (.CLK(clk_L0_B2), .D([2517]), .Q([554]), .Q_N([3000]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5140 (.CLK(clk_L0_B2), .D([2522]), .Q([552]), .Q_N([3001]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5141 (.CLK(clk_L0_B2), .D([2525]), .Q([453]), .Q_N([3002]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5142 (.CLK(clk_L0_B2), .D([2528]), .Q([454]), .Q_N([3003]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5143 (.CLK(clk_L0_B2), .D([2531]), .Q([2021]), .Q_N([3004]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5144 (.CLK(clk_L0_B2), .D([2534]), .Q([2014]), .Q_N([3005]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5145 (.CLK(clk_L0_B2), .D([2538]), .Q([2138]), .Q_N([3006]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5146 (.CLK(clk_L0_B2), .D([2543]), .Q([511]), .Q_N([3007]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5151 (.CLK(clk_L0_B2), .D([2552]), .Q([1523]), .Q_N([3008]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5152 (.CLK(clk_L0_B2), .D([2555]), .Q([1555]), .Q_N([3009]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5153 (.CLK(clk_L0_B2), .D([2566]), .Q([544]), .Q_N([3010]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5154 (.CLK(clk_L0_B2), .D([2568]), .Q([539]), .Q_N([3011]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5155 (.CLK(clk_L0_B4), .D([2574]), .Q([546]), .Q_N([3012]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5156 (.CLK(clk_L0_B4), .D([2578]), .Q([1886]), .Q_N([2197]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5157 (.CLK(clk_L0_B4), .D([2584]), .Q([1543]), .Q_N([3013]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5158 (.CLK(clk_L0_B4), .D([2587]), .Q([1525]), .Q_N([3014]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5159 (.CLK(clk_L0_B4), .D([2591]), .Q([1196]), .Q_N([562]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5160 (.CLK(clk_L0_B4), .D([2597]), .Q([1193]), .Q_N([3015]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5161 (.CLK(clk_L0_B4), .D([2606]), .Q([2175]), .Q_N([3016]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5166 (.CLK(clk_L0_B4), .D([2629]), .Q([481]), .Q_N([3017]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5167 (.CLK(clk_L0_B4), .D([2667]), .Q([675]), .Q_N([3018]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5168 (.CLK(clk_L0_B4), .D([2685]), .Q([721]), .Q_N([3019]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5169 (.CLK(clk_L0_B4), .D([141]), .Q([138]), .Q_N([3020]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5170 (.CLK(clk_L0_B4), .D([166]), .Q([142]), .Q_N([3021]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5171 (.CLK(clk_L0_B4), .D([188]), .Q([167]), .Q_N([3022]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5172 (.CLK(clk_L0_B4), .D([210]), .Q([189]), .Q_N([3023]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5173 (.CLK(clk_L0_B4), .D([231]), .Q([211]), .Q_N([3024]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5174 (.CLK(clk_L0_B4), .D([252]), .Q([232]), .Q_N([3025]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5175 (.CLK(clk_L0_B5), .D([278]), .Q([253]), .Q_N([3026]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5176 (.CLK(clk_L0_B6), .D([302]), .Q([279]), .Q_N([3027]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5177 (.CLK(clk_L0_B6), .D([326]), .Q([303]), .Q_N([3028]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5178 (.CLK(clk_L0_B6), .D([348]), .Q([327]), .Q_N([3029]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5179 (.CLK(clk_L0_B6), .D([372]), .Q([349]), .Q_N([3030]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5180 (.CLK(clk_L0_B6), .D([395]), .Q([373]), .Q_N([3031]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5181 (.CLK(clk_L0_B6), .D([416]), .Q([396]), .Q_N([3032]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5182 (.CLK(clk_L0_B6), .D([437]), .Q([417]), .Q_N([3033]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5183 (.CLK(clk_L0_B6), .D([1998]), .Q([1995]), .Q_N([2672]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5189 (.CLK(clk_L0_B6), .D([256]), .Q([2214]), .Q_N([3034]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5190 (.CLK(clk_L0_B5), .D([281]), .Q([2231]), .Q_N([3035]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5191 (.CLK(clk_L0_B5), .D([305]), .Q([2250]), .Q_N([3036]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5192 (.CLK(clk_L0_B5), .D([329]), .Q([2269]), .Q_N([3037]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5193 (.CLK(clk_L0_B5), .D([352]), .Q([2294]), .Q_N([3038]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5194 (.CLK(clk_L0_B5), .D([375]), .Q([2310]), .Q_N([3039]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5195 (.CLK(clk_L0_B5), .D([398]), .Q([2329]), .Q_N([3040]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5196 (.CLK(clk_L0_B5), .D([419]), .Q([2347]), .Q_N([3041]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5197 (.CLK(clk_L0_B5), .D([442]), .Q([438]), .Q_N([1238]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5198 (.CLK(clk_L0_B5), .D([447]), .Q([443]), .Q_N([1232]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5199 (.CLK(clk_L0_B5), .D([452]), .Q([448]), .Q_N([2148]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5200 (.CLK(clk_L0_B5), .D([2008]), .Q([2000]), .Q_N([3042]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5201 (.CLK(clk_L0_B5), .D([480]), .Q([474]), .Q_N([3043]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5202 (.CLK(clk_L0_B5), .D([507]), .Q([2121]), .Q_N([1249]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5203 (.CLK(clk_L0_B5), .D([2030]), .Q([2009]), .Q_N([2467]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5204 (.CLK(clk_L0_B5), .D([538]), .Q([531]), .Q_N([1235]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5205 (.CLK(clk_L0_B6), .D([582]), .Q([577]), .Q_N([1230]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5206 (.CLK(clk_L0_B6), .D([586]), .Q([583]), .Q_N([3044]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5207 (.CLK(clk_L0_B6), .D([704]), .Q([678]), .Q_N([3045]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5208 (.CLK(clk_L0_B6), .D([735]), .Q([724]), .Q_N([3046]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5209 (.CLK(clk_L0_B6), .D([765]), .Q([753]), .Q_N([3047]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5210 (.CLK(clk_L0_B6), .D([794]), .Q([152]), .Q_N([3048]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5211 (.CLK(clk_L0_B6), .D([823]), .Q([175]), .Q_N([3049]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5212 (.CLK(clk_L0_B7), .D([852]), .Q([194]), .Q_N([3050]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5213 (.CLK(clk_L0_B7), .D([881]), .Q([218]), .Q_N([3051]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5214 (.CLK(clk_L0_B7), .D([908]), .Q([239]), .Q_N([3052]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5215 (.CLK(clk_L0_B7), .D([2133]), .Q([3053]), .Q_N([2196]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5216 (.CLK(clk_L0_B7), .D([921]), .Q([258]), .Q_N([3054]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5217 (.CLK(clk_L0_B7), .D([932]), .Q([283]), .Q_N([3055]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5218 (.CLK(clk_L0_B7), .D([943]), .Q([307]), .Q_N([3056]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5219 (.CLK(clk_L0_B7), .D([954]), .Q([331]), .Q_N([3057]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5220 (.CLK(clk_L0_B7), .D([965]), .Q([355]), .Q_N([3058]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5221 (.CLK(clk_L0_B7), .D([976]), .Q([378]), .Q_N([3059]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5222 (.CLK(clk_L0_B7), .D([989]), .Q([400]), .Q_N([3060]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5223 (.CLK(clk_L0_B7), .D([1000]), .Q([421]), .Q_N([3061]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5224 (.CLK(clk_L0_B7), .D([1008]), .Q([1006]), .Q_N([3062]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5225 (.CLK(clk_L0_B7), .D([1012]), .Q([1010]), .Q_N([3063]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5226 (.CLK(clk_L0_B7), .D([1017]), .Q([1013]), .Q_N([3064]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5227 (.CLK(clk_L0_B7), .D([1021]), .Q([1019]), .Q_N([3065]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5228 (.CLK(clk_L0_B8), .D([1025]), .Q([1023]), .Q_N([3066]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5229 (.CLK(clk_L0_B8), .D([1030]), .Q([1026]), .Q_N([3067]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5230 (.CLK(clk_L0_B8), .D([1035]), .Q([1031]), .Q_N([3068]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5231 (.CLK(clk_L0_B8), .D([1039]), .Q([1036]), .Q_N([3069]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5232 (.CLK(clk_L0_B8), .D([1218]), .Q([1216]), .Q_N([2158]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5233 (.CLK(clk_L0_B8), .D([1291]), .Q([1288]), .Q_N([2150]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5234 (.CLK(clk_L0_B8), .D([1318]), .Q([1316]), .Q_N([2159]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5235 (.CLK(clk_L0_B8), .D([1348]), .Q([1346]), .Q_N([2152]), .RESET_B([2694]), .SET_B([3]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5236 (.CLK(clk_L0_B8), .D([1370]), .Q([1368]), .Q_N([2155]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5237 (.CLK(clk_L0_B8), .D([1385]), .Q([1383]), .Q_N([2149]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8804 (.CLK(clk_L0_B8), .D([1409]), .Q([1386]), .Q_N([3070]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8805 (.CLK(clk_L0_B8), .D([1421]), .Q([1410]), .Q_N([3071]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8806 (.CLK(clk_L0_B8), .D([1444]), .Q([2147]), .Q_N([3072]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8807 (.CLK(clk_L0_B8), .D([1452]), .Q([1449]), .Q_N([3073]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8808 (.CLK(clk_L0_B8), .D([1472]), .Q([1453]), .Q_N([3074]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8809 (.CLK(clk_L0_B8), .D([1490]), .Q([1488]), .Q_N([3075]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8810 (.CLK(clk_L0_B9), .D([1503]), .Q([1491]), .Q_N([3076]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8811 (.CLK(clk_L0_B9), .D([1512]), .Q([1504]), .Q_N([3077]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7456 (.CLK(clk_L0_B9), .D([1653]), .Q([1513]), .Q_N([3078]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7679 (.CLK(clk_L0_B9), .D([1922]), .Q([234]), .Q_N([3079]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7680 (.CLK(clk_L0_B9), .D([1926]), .Q([1923]), .Q_N([2199]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7681 (.CLK(clk_L0_B9), .D([1932]), .Q([516]), .Q_N([3080]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7682 (.CLK(clk_L0_B9), .D([1936]), .Q([286]), .Q_N([3081]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7683 (.CLK(clk_L0_B9), .D([1940]), .Q([518]), .Q_N([3082]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7684 (.CLK(clk_L0_B9), .D([1944]), .Q([145]), .Q_N([3083]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7685 (.CLK(clk_L0_B9), .D([1950]), .Q([169]), .Q_N([3084]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7686 (.CLK(clk_L0_B9), .D([1956]), .Q([191]), .Q_N([3085]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7687 (.CLK(clk_L0_B9), .D([1962]), .Q([213]), .Q_N([3086]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7689 (.CLK(clk_L0_B9), .D([1966]), .Q([1963]), .Q_N([3087]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7690 (.CLK(clk_L0_B9), .D([1982]), .Q([550]), .Q_N([2279]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__clkbuf_4 T0Y0__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B10));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R0_INV_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y0__R1_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B45));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R1_INV_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R2_INV_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R2_INV_1 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y0__R3_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B5));
  sky130_fd_sc_hd__clkbuf_4 T0Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1081));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R0_INV_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y10__R1_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1117));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R1_INV_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R2_INV_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R2_INV_1 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1153));
  sky130_fd_sc_hd__clkbuf_4 T0Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1189));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R0_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1225));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R1_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R2_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R2_INV_1 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y11__R3_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1261));
  sky130_fd_sc_hd__clkbuf_4 T0Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1297));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R0_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1333));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R1_INV_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R2_INV_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R2_INV_1 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1369));
  sky130_fd_sc_hd__clkbuf_4 T0Y13__R0_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1405));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R0_INV_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1441));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R1_INV_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R2_INV_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R2_INV_1 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1477));
  sky130_fd_sc_hd__clkbuf_4 T0Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1513));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R0_INV_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y14__R1_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B3));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R1_INV_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R2_INV_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R2_INV_1 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y14__R3_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B99));
  sky130_fd_sc_hd__clkbuf_4 T0Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1620));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R0_INV_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1656));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R1_INV_0 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R2_INV_0 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R2_INV_1 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y15__R3_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1692));
  sky130_fd_sc_hd__clkbuf_4 T0Y16__R0_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B108));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R0_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1764));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R1_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R2_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R2_INV_1 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1800));
  sky130_fd_sc_hd__clkbuf_4 T0Y17__R0_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1836));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R0_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y17__R1_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B117));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R1_INV_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R2_INV_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R2_INV_1 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1908));
  sky130_fd_sc_hd__clkbuf_4 T0Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1944));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R0_INV_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y18__R1_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1980));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R1_INV_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R2_INV_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R2_INV_1 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y18__R3_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B126));
  sky130_fd_sc_hd__clkbuf_4 T0Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2052));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R0_INV_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2088));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R1_INV_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R2_INV_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R2_INV_1 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y19__R3_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2124));
  sky130_fd_sc_hd__clkbuf_4 T0Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B115));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R0_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B150));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R1_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R2_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R2_INV_1 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B185));
  sky130_fd_sc_hd__clkbuf_4 T0Y20__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B135));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R0_INV_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2196));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R1_INV_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R2_INV_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R2_INV_1 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2232));
  sky130_fd_sc_hd__clkbuf_4 T0Y21__R0_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2268));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R0_INV_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y21__R1_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B9));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R1_INV_0 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R2_INV_0 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R2_INV_1 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2340));
  sky130_fd_sc_hd__clkbuf_4 T0Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2376));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R0_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y22__R1_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2412));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R1_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R2_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R2_INV_1 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y22__R3_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B153));
  sky130_fd_sc_hd__clkbuf_4 T0Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2484));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R0_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2520));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R1_INV_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R2_INV_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R2_INV_1 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y23__R3_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2556));
  sky130_fd_sc_hd__clkbuf_4 T0Y24__R0_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B162));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R0_INV_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2628));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R1_INV_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R2_INV_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R2_INV_1 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2664));
  sky130_fd_sc_hd__clkbuf_4 T0Y25__R0_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2700));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R0_INV_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y25__R1_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B171));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R1_INV_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R2_INV_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R2_INV_1 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2772));
  sky130_fd_sc_hd__clkbuf_4 T0Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2808));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R0_INV_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y26__R1_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2844));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R1_INV_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R2_INV_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R2_INV_1 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y26__R3_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B180));
  sky130_fd_sc_hd__clkbuf_4 T0Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2916));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R0_INV_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2952));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R1_INV_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R2_INV_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R2_INV_1 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y27__R3_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2988));
  sky130_fd_sc_hd__clkbuf_4 T0Y28__R0_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B189));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R0_INV_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3060));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R1_INV_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R2_INV_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R2_INV_1 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3096));
  sky130_fd_sc_hd__clkbuf_4 T0Y29__R0_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3132));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R0_INV_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y29__R1_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B198));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R1_INV_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R2_INV_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R2_INV_1 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3204));
  sky130_fd_sc_hd__clkbuf_4 T0Y2__R0_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B220));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R0_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y2__R1_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B255));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R1_INV_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R2_INV_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R2_INV_1 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B291));
  sky130_fd_sc_hd__clkbuf_4 T0Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3240));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R0_INV_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y30__R1_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3276));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R1_INV_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R2_INV_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R2_INV_1 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y30__R3_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B207));
  sky130_fd_sc_hd__clkbuf_4 T0Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3348));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R0_INV_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3384));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R1_INV_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R2_INV_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R2_INV_1 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y31__R3_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3420));
  sky130_fd_sc_hd__clkbuf_4 T0Y32__R0_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B216));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R0_INV_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3492));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R1_INV_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R2_INV_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R2_INV_1 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3528));
  sky130_fd_sc_hd__clkbuf_4 T0Y33__R0_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3564));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R0_INV_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y33__R1_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B225));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R1_INV_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R2_INV_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R2_INV_1 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3636));
  sky130_fd_sc_hd__clkbuf_4 T0Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3672));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R0_INV_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y34__R1_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3708));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R1_INV_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R2_INV_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R2_INV_1 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y34__R3_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B234));
  sky130_fd_sc_hd__clkbuf_4 T0Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3780));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R0_INV_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3816));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R1_INV_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R2_INV_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R2_INV_1 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y35__R3_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3852));
  sky130_fd_sc_hd__clkbuf_4 T0Y36__R0_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B243));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R0_INV_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3924));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R1_INV_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R2_INV_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R2_INV_1 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3960));
  sky130_fd_sc_hd__clkbuf_4 T0Y37__R0_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3996));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R0_INV_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y37__R1_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B252));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R1_INV_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R2_INV_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R2_INV_1 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4068));
  sky130_fd_sc_hd__clkbuf_4 T0Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4104));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R0_INV_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y38__R1_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4140));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R1_INV_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R2_INV_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R2_INV_1 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y38__R3_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B261));
  sky130_fd_sc_hd__clkbuf_4 T0Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4212));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R0_INV_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4248));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R1_INV_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R2_INV_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R2_INV_1 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y39__R3_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4284));
  sky130_fd_sc_hd__clkbuf_4 T0Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B326));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R0_INV_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B361));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R1_INV_0 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R2_INV_0 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R2_INV_1 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y3__R3_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B397));
  sky130_fd_sc_hd__clkbuf_4 T0Y40__R0_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B270));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R0_INV_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4356));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R1_INV_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R2_INV_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R2_INV_1 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4392));
  sky130_fd_sc_hd__clkbuf_4 T0Y41__R0_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4428));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R0_INV_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y41__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B279));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R1_INV_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R2_INV_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R2_INV_1 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4500));
  sky130_fd_sc_hd__clkbuf_4 T0Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4536));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R0_INV_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y42__R1_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4572));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R1_INV_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R2_INV_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R2_INV_1 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y42__R3_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B18));
  sky130_fd_sc_hd__clkbuf_4 T0Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4644));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R0_INV_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4680));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R1_INV_0 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R2_INV_0 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R2_INV_1 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y43__R3_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4716));
  sky130_fd_sc_hd__clkbuf_4 T0Y44__R0_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B297));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R0_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4788));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R1_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R2_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R2_INV_1 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4824));
  sky130_fd_sc_hd__clkbuf_4 T0Y45__R0_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4860));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R0_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y45__R1_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B306));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R1_INV_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R2_INV_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R2_INV_1 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4932));
  sky130_fd_sc_hd__clkbuf_4 T0Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4968));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R0_INV_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y46__R1_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5004));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R1_INV_0 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R2_INV_0 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R2_INV_1 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y46__R3_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B315));
  sky130_fd_sc_hd__clkbuf_4 T0Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5076));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R0_INV_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5112));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R1_INV_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R2_INV_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R2_INV_1 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y47__R3_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5148));
  sky130_fd_sc_hd__clkbuf_4 T0Y48__R0_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B324));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R0_INV_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5220));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R1_INV_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R2_INV_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R2_INV_1 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5256));
  sky130_fd_sc_hd__clkbuf_4 T0Y49__R0_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5292));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R0_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y49__R1_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B333));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R1_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R2_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R2_INV_1 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5364));
  sky130_fd_sc_hd__clkbuf_4 T0Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B433));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R0_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B469));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R1_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R2_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R2_INV_1 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B505));
  sky130_fd_sc_hd__clkbuf_4 T0Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5400));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R0_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y50__R1_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5436));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R1_INV_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R2_INV_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R2_INV_1 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y50__R3_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B342));
  sky130_fd_sc_hd__clkbuf_4 T0Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5508));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R0_INV_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5544));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R1_INV_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R2_INV_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R2_INV_1 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y51__R3_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5580));
  sky130_fd_sc_hd__clkbuf_4 T0Y52__R0_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B351));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R0_INV_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5652));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R1_INV_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R2_INV_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R2_INV_1 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5688));
  sky130_fd_sc_hd__clkbuf_4 T0Y53__R0_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5724));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R0_INV_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y53__R1_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B360));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R1_INV_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R2_INV_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R2_INV_1 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5796));
  sky130_fd_sc_hd__clkbuf_4 T0Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5832));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R0_INV_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y54__R1_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5868));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R1_INV_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R2_INV_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R2_INV_1 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y54__R3_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B369));
  sky130_fd_sc_hd__clkbuf_4 T0Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5940));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R0_INV_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5976));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R1_INV_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R2_INV_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R2_INV_1 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y55__R3_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6012));
  sky130_fd_sc_hd__clkbuf_4 T0Y56__R0_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B378));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R0_INV_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6084));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R1_INV_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R2_INV_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R2_INV_1 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6120));
  sky130_fd_sc_hd__clkbuf_4 T0Y57__R0_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6156));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R0_INV_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y57__R1_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B387));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R1_INV_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R2_INV_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R2_INV_1 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6228));
  sky130_fd_sc_hd__clkbuf_4 T0Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6264));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R0_INV_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y58__R1_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6300));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R1_INV_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R2_INV_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R2_INV_1 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y58__R3_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B396));
  sky130_fd_sc_hd__clkbuf_4 T0Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6372));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R0_INV_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6408));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R1_INV_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R2_INV_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R2_INV_1 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y59__R3_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6444));
  sky130_fd_sc_hd__clkbuf_4 T0Y5__R0_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B541));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R0_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B577));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R1_INV_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R2_INV_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R2_INV_1 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B613));
  sky130_fd_sc_hd__clkbuf_4 T0Y60__R0_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B405));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R0_INV_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6516));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R1_INV_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R2_INV_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R2_INV_1 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6552));
  sky130_fd_sc_hd__clkbuf_4 T0Y61__R0_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6588));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R0_INV_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y61__R1_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B414));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R1_INV_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R2_INV_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R2_INV_1 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6660));
  sky130_fd_sc_hd__clkbuf_4 T0Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6696));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R0_INV_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y62__R1_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6732));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R1_INV_0 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R2_INV_0 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R2_INV_1 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y62__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B423));
  sky130_fd_sc_hd__clkbuf_4 T0Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6804));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R0_INV_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6840));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R1_INV_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R2_INV_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R2_INV_1 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y63__R3_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6876));
  sky130_fd_sc_hd__clkbuf_4 T0Y64__R0_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B27));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R0_INV_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6948));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R1_INV_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R2_INV_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R2_INV_1 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6984));
  sky130_fd_sc_hd__clkbuf_4 T0Y65__R0_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7020));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R0_INV_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y65__R1_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B441));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R1_INV_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R2_INV_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R2_INV_1 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7092));
  sky130_fd_sc_hd__clkbuf_4 T0Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7128));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R0_INV_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y66__R1_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7164));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R1_INV_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R2_INV_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R2_INV_1 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y66__R3_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B450));
  sky130_fd_sc_hd__clkbuf_4 T0Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7236));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R0_INV_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7272));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R1_INV_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R2_INV_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R2_INV_1 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y67__R3_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7308));
  sky130_fd_sc_hd__clkbuf_4 T0Y68__R0_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B459));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R0_INV_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7380));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R1_INV_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R2_INV_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R2_INV_1 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7416));
  sky130_fd_sc_hd__clkbuf_4 T0Y69__R0_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7452));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R0_INV_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y69__R1_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B468));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R1_INV_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R2_INV_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R2_INV_1 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7524));
  sky130_fd_sc_hd__clkbuf_4 T0Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B649));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R0_INV_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y6__R1_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B685));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R1_INV_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R2_INV_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R2_INV_1 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B721));
  sky130_fd_sc_hd__clkbuf_4 T0Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7560));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R0_INV_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y70__R1_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7596));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R1_INV_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R2_INV_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R2_INV_1 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y70__R3_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B477));
  sky130_fd_sc_hd__clkbuf_4 T0Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7668));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R0_INV_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7704));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R1_INV_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R2_INV_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R2_INV_1 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y71__R3_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7740));
  sky130_fd_sc_hd__clkbuf_4 T0Y72__R0_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B486));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R0_INV_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7812));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R1_INV_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R2_INV_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R2_INV_1 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7848));
  sky130_fd_sc_hd__clkbuf_4 T0Y73__R0_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7884));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R0_INV_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y73__R1_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B495));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R1_INV_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R2_INV_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R2_INV_1 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7956));
  sky130_fd_sc_hd__clkbuf_4 T0Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7992));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R0_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y74__R1_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8028));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R1_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R2_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R2_INV_1 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y74__R3_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B504));
  sky130_fd_sc_hd__clkbuf_4 T0Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8100));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R0_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8136));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R1_INV_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R2_INV_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R2_INV_1 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y75__R3_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8172));
  sky130_fd_sc_hd__clkbuf_4 T0Y76__R0_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B513));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R0_INV_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8244));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R1_INV_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R2_INV_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R2_INV_1 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8280));
  sky130_fd_sc_hd__clkbuf_4 T0Y77__R0_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8316));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R0_INV_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y77__R1_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B522));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R1_INV_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R2_INV_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R2_INV_1 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8388));
  sky130_fd_sc_hd__clkbuf_4 T0Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8424));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R0_INV_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y78__R1_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8460));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R1_INV_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R2_INV_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R2_INV_1 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y78__R3_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B531));
  sky130_fd_sc_hd__clkbuf_4 T0Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8532));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R0_INV_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8568));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R1_INV_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R2_INV_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R2_INV_1 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y79__R3_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8604));
  sky130_fd_sc_hd__clkbuf_4 T0Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B757));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R0_INV_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B793));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R1_INV_0 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R2_INV_0 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R2_INV_1 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y7__R3_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B829));
  sky130_fd_sc_hd__clkbuf_4 T0Y80__R0_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B540));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R0_INV_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8676));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R1_INV_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R2_INV_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R2_INV_1 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8712));
  sky130_fd_sc_hd__clkbuf_4 T0Y81__R0_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8748));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R0_INV_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y81__R1_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B549));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R1_INV_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R2_INV_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R2_INV_1 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8820));
  sky130_fd_sc_hd__clkbuf_4 T0Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8856));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R0_INV_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y82__R1_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8892));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R1_INV_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R2_INV_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R2_INV_1 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y82__R3_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B558));
  sky130_fd_sc_hd__clkbuf_4 T0Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8964));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R0_INV_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9000));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R1_INV_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R2_INV_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R2_INV_1 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y83__R3_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9036));
  sky130_fd_sc_hd__clkbuf_4 T0Y84__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B567));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R0_INV_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9108));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R1_INV_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R2_INV_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R2_INV_1 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9144));
  sky130_fd_sc_hd__clkbuf_4 T0Y85__R0_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9180));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R0_INV_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y85__R1_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B36));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R1_INV_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R2_INV_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R2_INV_1 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9252));
  sky130_fd_sc_hd__clkbuf_4 T0Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9288));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R0_INV_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y86__R1_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9324));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R1_INV_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R2_INV_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R2_INV_1 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y86__R3_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B585));
  sky130_fd_sc_hd__clkbuf_4 T0Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9396));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R0_INV_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9432));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R1_INV_0 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R2_INV_0 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R2_INV_1 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y87__R3_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9468));
  sky130_fd_sc_hd__clkbuf_4 T0Y88__R0_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B594));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R0_INV_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9540));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R1_INV_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R2_INV_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R2_INV_1 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9576));
  sky130_fd_sc_hd__clkbuf_4 T0Y89__R0_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9612));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R0_INV_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y89__R1_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B603));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R1_INV_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R2_INV_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R2_INV_1 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9684));
  sky130_fd_sc_hd__clkbuf_4 T0Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B865));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R0_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B901));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R1_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R2_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R2_INV_1 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B937));
  sky130_fd_sc_hd__clkbuf_4 T0Y9__R0_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B973));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R0_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1009));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R1_INV_0 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R2_INV_0 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R2_INV_1 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1045));
  sky130_fd_sc_hd__clkbuf_4 T10Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B20));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R0_INV_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B55));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R1_INV_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R2_INV_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R2_INV_1 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B90));
  sky130_fd_sc_hd__clkbuf_4 T10Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1091));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R0_INV_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1127));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R1_INV_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R2_INV_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R2_INV_1 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1163));
  sky130_fd_sc_hd__clkbuf_4 T10Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1199));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R0_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1235));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R1_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R2_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R2_INV_1 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1271));
  sky130_fd_sc_hd__clkbuf_4 T10Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1307));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R0_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1343));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R1_INV_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R2_INV_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R2_INV_1 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1379));
  sky130_fd_sc_hd__clkbuf_4 T10Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1415));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R0_INV_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1451));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R1_INV_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R2_INV_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R2_INV_1 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1487));
  sky130_fd_sc_hd__clkbuf_4 T10Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1523));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R0_INV_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1558));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R1_INV_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R2_INV_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R2_INV_1 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1594));
  sky130_fd_sc_hd__clkbuf_4 T10Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1630));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R0_INV_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1666));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R1_INV_0 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R2_INV_0 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R2_INV_1 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1702));
  sky130_fd_sc_hd__clkbuf_4 T10Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1738));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R0_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1774));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R1_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R2_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R2_INV_1 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1810));
  sky130_fd_sc_hd__clkbuf_4 T10Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1846));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R0_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1882));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R1_INV_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R2_INV_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R2_INV_1 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1918));
  sky130_fd_sc_hd__clkbuf_4 T10Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1954));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R0_INV_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1990));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R1_INV_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R2_INV_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R2_INV_1 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2026));
  sky130_fd_sc_hd__clkbuf_4 T10Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2062));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R0_INV_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2098));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R1_INV_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R2_INV_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R2_INV_1 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2134));
  sky130_fd_sc_hd__clkbuf_4 T10Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B125));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R0_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y1__R1_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B10));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R1_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R2_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R2_INV_1 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B195));
  sky130_fd_sc_hd__clkbuf_4 T10Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2170));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R0_INV_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2206));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R1_INV_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R2_INV_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R2_INV_1 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2242));
  sky130_fd_sc_hd__clkbuf_4 T10Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2278));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R0_INV_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2314));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R1_INV_0 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R2_INV_0 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R2_INV_1 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2350));
  sky130_fd_sc_hd__clkbuf_4 T10Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2386));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R0_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2422));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R1_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R2_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R2_INV_1 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2458));
  sky130_fd_sc_hd__clkbuf_4 T10Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2494));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R0_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2530));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R1_INV_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R2_INV_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R2_INV_1 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2566));
  sky130_fd_sc_hd__clkbuf_4 T10Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2602));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R0_INV_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2638));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R1_INV_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R2_INV_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R2_INV_1 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2674));
  sky130_fd_sc_hd__clkbuf_4 T10Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2710));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R0_INV_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2746));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R1_INV_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R2_INV_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R2_INV_1 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2782));
  sky130_fd_sc_hd__clkbuf_4 T10Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2818));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R0_INV_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2854));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R1_INV_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R2_INV_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R2_INV_1 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2890));
  sky130_fd_sc_hd__clkbuf_4 T10Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2926));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R0_INV_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2962));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R1_INV_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R2_INV_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R2_INV_1 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2998));
  sky130_fd_sc_hd__clkbuf_4 T10Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3034));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R0_INV_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3070));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R1_INV_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R2_INV_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R2_INV_1 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3106));
  sky130_fd_sc_hd__clkbuf_4 T10Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3142));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R0_INV_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3178));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R1_INV_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R2_INV_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R2_INV_1 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3214));
  sky130_fd_sc_hd__clkbuf_4 T10Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B230));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R0_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B265));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R1_INV_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R2_INV_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R2_INV_1 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B301));
  sky130_fd_sc_hd__clkbuf_4 T10Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3250));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R0_INV_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3286));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R1_INV_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R2_INV_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R2_INV_1 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3322));
  sky130_fd_sc_hd__clkbuf_4 T10Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3358));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R0_INV_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3394));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R1_INV_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R2_INV_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R2_INV_1 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3430));
  sky130_fd_sc_hd__clkbuf_4 T10Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3466));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R0_INV_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3502));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R1_INV_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R2_INV_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R2_INV_1 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3538));
  sky130_fd_sc_hd__clkbuf_4 T10Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3574));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R0_INV_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3610));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R1_INV_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R2_INV_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R2_INV_1 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3646));
  sky130_fd_sc_hd__clkbuf_4 T10Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3682));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R0_INV_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3718));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R1_INV_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R2_INV_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R2_INV_1 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3754));
  sky130_fd_sc_hd__clkbuf_4 T10Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3790));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R0_INV_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3826));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R1_INV_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R2_INV_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R2_INV_1 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3862));
  sky130_fd_sc_hd__clkbuf_4 T10Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3898));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R0_INV_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3934));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R1_INV_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R2_INV_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R2_INV_1 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3970));
  sky130_fd_sc_hd__clkbuf_4 T10Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4006));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R0_INV_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4042));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R1_INV_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R2_INV_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R2_INV_1 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4078));
  sky130_fd_sc_hd__clkbuf_4 T10Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4114));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R0_INV_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4150));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R1_INV_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R2_INV_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R2_INV_1 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4186));
  sky130_fd_sc_hd__clkbuf_4 T10Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4222));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R0_INV_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4258));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R1_INV_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R2_INV_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R2_INV_1 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4294));
  sky130_fd_sc_hd__clkbuf_4 T10Y3__R0_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B21));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R0_INV_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B371));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R1_INV_0 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R2_INV_0 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R2_INV_1 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B407));
  sky130_fd_sc_hd__clkbuf_4 T10Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4330));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R0_INV_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4366));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R1_INV_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R2_INV_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R2_INV_1 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4402));
  sky130_fd_sc_hd__clkbuf_4 T10Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4438));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R0_INV_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4474));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R1_INV_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R2_INV_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R2_INV_1 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4510));
  sky130_fd_sc_hd__clkbuf_4 T10Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4546));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R0_INV_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4582));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R1_INV_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R2_INV_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R2_INV_1 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4618));
  sky130_fd_sc_hd__clkbuf_4 T10Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4654));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R0_INV_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4690));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R1_INV_0 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R2_INV_0 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R2_INV_1 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4726));
  sky130_fd_sc_hd__clkbuf_4 T10Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4762));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R0_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4798));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R1_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R2_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R2_INV_1 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4834));
  sky130_fd_sc_hd__clkbuf_4 T10Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4870));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R0_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4906));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R1_INV_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R2_INV_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R2_INV_1 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4942));
  sky130_fd_sc_hd__clkbuf_4 T10Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4978));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R0_INV_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5014));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R1_INV_0 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R2_INV_0 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R2_INV_1 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5050));
  sky130_fd_sc_hd__clkbuf_4 T10Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5086));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R0_INV_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5122));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R1_INV_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R2_INV_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R2_INV_1 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5158));
  sky130_fd_sc_hd__clkbuf_4 T10Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5194));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R0_INV_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5230));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R1_INV_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R2_INV_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R2_INV_1 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5266));
  sky130_fd_sc_hd__clkbuf_4 T10Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5302));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R0_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5338));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R1_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R2_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R2_INV_1 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5374));
  sky130_fd_sc_hd__clkbuf_4 T10Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B443));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R0_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B479));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R1_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R2_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R2_INV_1 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B515));
  sky130_fd_sc_hd__clkbuf_4 T10Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5410));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R0_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5446));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R1_INV_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R2_INV_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R2_INV_1 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5482));
  sky130_fd_sc_hd__clkbuf_4 T10Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5518));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R0_INV_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5554));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R1_INV_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R2_INV_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R2_INV_1 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5590));
  sky130_fd_sc_hd__clkbuf_4 T10Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5626));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R0_INV_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5662));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R1_INV_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R2_INV_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R2_INV_1 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5698));
  sky130_fd_sc_hd__clkbuf_4 T10Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5734));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R0_INV_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5770));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R1_INV_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R2_INV_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R2_INV_1 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5806));
  sky130_fd_sc_hd__clkbuf_4 T10Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5842));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R0_INV_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5878));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R1_INV_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R2_INV_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R2_INV_1 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5914));
  sky130_fd_sc_hd__clkbuf_4 T10Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5950));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R0_INV_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5986));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R1_INV_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R2_INV_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R2_INV_1 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6022));
  sky130_fd_sc_hd__clkbuf_4 T10Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6058));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R0_INV_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6094));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R1_INV_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R2_INV_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R2_INV_1 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6130));
  sky130_fd_sc_hd__clkbuf_4 T10Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6166));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R0_INV_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6202));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R1_INV_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R2_INV_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R2_INV_1 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6238));
  sky130_fd_sc_hd__clkbuf_4 T10Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6274));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R0_INV_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6310));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R1_INV_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R2_INV_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R2_INV_1 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6346));
  sky130_fd_sc_hd__clkbuf_4 T10Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6382));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R0_INV_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6418));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R1_INV_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R2_INV_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R2_INV_1 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6454));
  sky130_fd_sc_hd__clkbuf_4 T10Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B551));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R0_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B587));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R1_INV_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R2_INV_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R2_INV_1 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B623));
  sky130_fd_sc_hd__clkbuf_4 T10Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6490));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R0_INV_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6526));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R1_INV_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R2_INV_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R2_INV_1 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6562));
  sky130_fd_sc_hd__clkbuf_4 T10Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6598));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R0_INV_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6634));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R1_INV_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R2_INV_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R2_INV_1 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6670));
  sky130_fd_sc_hd__clkbuf_4 T10Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6706));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R0_INV_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6742));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R1_INV_0 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R2_INV_0 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R2_INV_1 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6778));
  sky130_fd_sc_hd__clkbuf_4 T10Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6814));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R0_INV_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6850));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R1_INV_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R2_INV_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R2_INV_1 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6886));
  sky130_fd_sc_hd__clkbuf_4 T10Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6922));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R0_INV_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6958));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R1_INV_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R2_INV_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R2_INV_1 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6994));
  sky130_fd_sc_hd__clkbuf_4 T10Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7030));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R0_INV_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7066));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R1_INV_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R2_INV_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R2_INV_1 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7102));
  sky130_fd_sc_hd__clkbuf_4 T10Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7138));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R0_INV_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7174));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R1_INV_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R2_INV_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R2_INV_1 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7210));
  sky130_fd_sc_hd__clkbuf_4 T10Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7246));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R0_INV_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7282));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R1_INV_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R2_INV_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R2_INV_1 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7318));
  sky130_fd_sc_hd__clkbuf_4 T10Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7354));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R0_INV_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7390));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R1_INV_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R2_INV_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R2_INV_1 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7426));
  sky130_fd_sc_hd__clkbuf_4 T10Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7462));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R0_INV_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7498));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R1_INV_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R2_INV_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R2_INV_1 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7534));
  sky130_fd_sc_hd__clkbuf_4 T10Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B659));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R0_INV_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B695));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R1_INV_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R2_INV_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R2_INV_1 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B731));
  sky130_fd_sc_hd__clkbuf_4 T10Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7570));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R0_INV_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7606));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R1_INV_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R2_INV_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R2_INV_1 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7642));
  sky130_fd_sc_hd__clkbuf_4 T10Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7678));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R0_INV_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7714));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R1_INV_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R2_INV_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R2_INV_1 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7750));
  sky130_fd_sc_hd__clkbuf_4 T10Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7786));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R0_INV_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7822));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R1_INV_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R2_INV_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R2_INV_1 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7858));
  sky130_fd_sc_hd__clkbuf_4 T10Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7894));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R0_INV_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7930));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R1_INV_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R2_INV_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R2_INV_1 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7966));
  sky130_fd_sc_hd__clkbuf_4 T10Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8002));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R0_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8038));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R1_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R2_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R2_INV_1 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8074));
  sky130_fd_sc_hd__clkbuf_4 T10Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8110));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R0_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8146));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R1_INV_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R2_INV_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R2_INV_1 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8182));
  sky130_fd_sc_hd__clkbuf_4 T10Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8218));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R0_INV_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8254));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R1_INV_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R2_INV_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R2_INV_1 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8290));
  sky130_fd_sc_hd__clkbuf_4 T10Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8326));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R0_INV_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8362));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R1_INV_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R2_INV_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R2_INV_1 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8398));
  sky130_fd_sc_hd__clkbuf_4 T10Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8434));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R0_INV_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8470));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R1_INV_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R2_INV_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R2_INV_1 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8506));
  sky130_fd_sc_hd__clkbuf_4 T10Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8542));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R0_INV_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8578));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R1_INV_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R2_INV_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R2_INV_1 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8614));
  sky130_fd_sc_hd__clkbuf_4 T10Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B767));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R0_INV_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B803));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R1_INV_0 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R2_INV_0 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R2_INV_1 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B839));
  sky130_fd_sc_hd__clkbuf_4 T10Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8650));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R0_INV_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8686));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R1_INV_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R2_INV_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R2_INV_1 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8722));
  sky130_fd_sc_hd__clkbuf_4 T10Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8758));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R0_INV_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8794));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R1_INV_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R2_INV_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R2_INV_1 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8830));
  sky130_fd_sc_hd__clkbuf_4 T10Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8866));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R0_INV_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8902));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R1_INV_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R2_INV_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R2_INV_1 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8938));
  sky130_fd_sc_hd__clkbuf_4 T10Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8974));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R0_INV_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9010));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R1_INV_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R2_INV_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R2_INV_1 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9046));
  sky130_fd_sc_hd__clkbuf_4 T10Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9082));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R0_INV_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9118));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R1_INV_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R2_INV_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R2_INV_1 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9154));
  sky130_fd_sc_hd__clkbuf_4 T10Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9190));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R0_INV_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9226));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R1_INV_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R2_INV_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R2_INV_1 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9262));
  sky130_fd_sc_hd__clkbuf_4 T10Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9298));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R0_INV_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9334));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R1_INV_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R2_INV_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R2_INV_1 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9370));
  sky130_fd_sc_hd__clkbuf_4 T10Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9406));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R0_INV_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9442));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R1_INV_0 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R2_INV_0 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R2_INV_1 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9478));
  sky130_fd_sc_hd__clkbuf_4 T10Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9514));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R0_INV_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9550));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R1_INV_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R2_INV_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R2_INV_1 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9586));
  sky130_fd_sc_hd__clkbuf_4 T10Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9622));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R0_INV_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9658));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R1_INV_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R2_INV_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R2_INV_1 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9694));
  sky130_fd_sc_hd__clkbuf_4 T10Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B875));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R0_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B911));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R1_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R2_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R2_INV_1 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B947));
  sky130_fd_sc_hd__clkbuf_4 T10Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B983));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R0_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1019));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R1_INV_0 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R2_INV_0 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R2_INV_1 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1055));
  sky130_fd_sc_hd__clkbuf_4 T11Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B21));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R0_INV_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B56));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R1_INV_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R2_INV_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R2_INV_1 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B91));
  sky130_fd_sc_hd__clkbuf_4 T11Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1092));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R0_INV_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1128));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R1_INV_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R2_INV_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R2_INV_1 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1164));
  sky130_fd_sc_hd__clkbuf_4 T11Y11__R0_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B75));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R0_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1236));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R1_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R2_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R2_INV_1 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1272));
  sky130_fd_sc_hd__clkbuf_4 T11Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1308));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R0_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y12__R1_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B84));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R1_INV_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R2_INV_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R2_INV_1 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1380));
  sky130_fd_sc_hd__clkbuf_4 T11Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1416));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R0_INV_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1452));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R1_INV_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R2_INV_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R2_INV_1 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y13__R3_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B93));
  sky130_fd_sc_hd__clkbuf_4 T11Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1524));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R0_INV_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1559));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R1_INV_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R2_INV_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R2_INV_1 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1595));
  sky130_fd_sc_hd__clkbuf_4 T11Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1631));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R0_INV_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1667));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R1_INV_0 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R2_INV_0 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R2_INV_1 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1703));
  sky130_fd_sc_hd__clkbuf_4 T11Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1739));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R0_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1775));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R1_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R2_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R2_INV_1 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1811));
  sky130_fd_sc_hd__clkbuf_4 T11Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1847));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R0_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1883));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R1_INV_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R2_INV_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R2_INV_1 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1919));
  sky130_fd_sc_hd__clkbuf_4 T11Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1955));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R0_INV_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1991));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R1_INV_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R2_INV_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R2_INV_1 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2027));
  sky130_fd_sc_hd__clkbuf_4 T11Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2063));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R0_INV_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2099));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R1_INV_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R2_INV_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R2_INV_1 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2135));
  sky130_fd_sc_hd__clkbuf_4 T11Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B126));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R0_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B161));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R1_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R2_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R2_INV_1 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B196));
  sky130_fd_sc_hd__clkbuf_4 T11Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2171));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R0_INV_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2207));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R1_INV_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R2_INV_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R2_INV_1 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2243));
  sky130_fd_sc_hd__clkbuf_4 T11Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2279));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R0_INV_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2315));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R1_INV_0 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R2_INV_0 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R2_INV_1 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2351));
  sky130_fd_sc_hd__clkbuf_4 T11Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2387));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R0_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2423));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R1_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R2_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R2_INV_1 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2459));
  sky130_fd_sc_hd__clkbuf_4 T11Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2495));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R0_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2531));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R1_INV_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R2_INV_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R2_INV_1 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2567));
  sky130_fd_sc_hd__clkbuf_4 T11Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2603));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R0_INV_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2639));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R1_INV_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R2_INV_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R2_INV_1 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2675));
  sky130_fd_sc_hd__clkbuf_4 T11Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2711));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R0_INV_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2747));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R1_INV_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R2_INV_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R2_INV_1 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2783));
  sky130_fd_sc_hd__clkbuf_4 T11Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2819));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R0_INV_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2855));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R1_INV_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R2_INV_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R2_INV_1 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2891));
  sky130_fd_sc_hd__clkbuf_4 T11Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2927));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R0_INV_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2963));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R1_INV_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R2_INV_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R2_INV_1 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2999));
  sky130_fd_sc_hd__clkbuf_4 T11Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3035));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R0_INV_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3071));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R1_INV_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R2_INV_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R2_INV_1 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3107));
  sky130_fd_sc_hd__clkbuf_4 T11Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3143));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R0_INV_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3179));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R1_INV_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R2_INV_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R2_INV_1 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3215));
  sky130_fd_sc_hd__clkbuf_4 T11Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B231));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R0_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B266));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R1_INV_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R2_INV_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R2_INV_1 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B302));
  sky130_fd_sc_hd__clkbuf_4 T11Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3251));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R0_INV_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3287));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R1_INV_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R2_INV_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R2_INV_1 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3323));
  sky130_fd_sc_hd__clkbuf_4 T11Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3359));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R0_INV_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3395));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R1_INV_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R2_INV_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R2_INV_1 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3431));
  sky130_fd_sc_hd__clkbuf_4 T11Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3467));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R0_INV_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3503));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R1_INV_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R2_INV_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R2_INV_1 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3539));
  sky130_fd_sc_hd__clkbuf_4 T11Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3575));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R0_INV_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3611));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R1_INV_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R2_INV_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R2_INV_1 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3647));
  sky130_fd_sc_hd__clkbuf_4 T11Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3683));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R0_INV_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3719));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R1_INV_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R2_INV_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R2_INV_1 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3755));
  sky130_fd_sc_hd__clkbuf_4 T11Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3791));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R0_INV_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3827));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R1_INV_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R2_INV_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R2_INV_1 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3863));
  sky130_fd_sc_hd__clkbuf_4 T11Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3899));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R0_INV_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3935));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R1_INV_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R2_INV_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R2_INV_1 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3971));
  sky130_fd_sc_hd__clkbuf_4 T11Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4007));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R0_INV_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4043));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R1_INV_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R2_INV_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R2_INV_1 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4079));
  sky130_fd_sc_hd__clkbuf_4 T11Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4115));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R0_INV_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4151));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R1_INV_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R2_INV_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R2_INV_1 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4187));
  sky130_fd_sc_hd__clkbuf_4 T11Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4223));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R0_INV_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4259));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R1_INV_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R2_INV_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R2_INV_1 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4295));
  sky130_fd_sc_hd__clkbuf_4 T11Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B337));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R0_INV_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B372));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R1_INV_0 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R2_INV_0 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R2_INV_1 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B408));
  sky130_fd_sc_hd__clkbuf_4 T11Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4331));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R0_INV_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4367));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R1_INV_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R2_INV_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R2_INV_1 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4403));
  sky130_fd_sc_hd__clkbuf_4 T11Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4439));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R0_INV_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4475));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R1_INV_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R2_INV_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R2_INV_1 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4511));
  sky130_fd_sc_hd__clkbuf_4 T11Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4547));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R0_INV_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4583));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R1_INV_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R2_INV_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R2_INV_1 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4619));
  sky130_fd_sc_hd__clkbuf_4 T11Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4655));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R0_INV_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4691));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R1_INV_0 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R2_INV_0 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R2_INV_1 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4727));
  sky130_fd_sc_hd__clkbuf_4 T11Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4763));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R0_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4799));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R1_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R2_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R2_INV_1 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4835));
  sky130_fd_sc_hd__clkbuf_4 T11Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4871));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R0_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4907));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R1_INV_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R2_INV_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R2_INV_1 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4943));
  sky130_fd_sc_hd__clkbuf_4 T11Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4979));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R0_INV_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5015));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R1_INV_0 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R2_INV_0 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R2_INV_1 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5051));
  sky130_fd_sc_hd__clkbuf_4 T11Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5087));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R0_INV_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5123));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R1_INV_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R2_INV_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R2_INV_1 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5159));
  sky130_fd_sc_hd__clkbuf_4 T11Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5195));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R0_INV_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5231));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R1_INV_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R2_INV_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R2_INV_1 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5267));
  sky130_fd_sc_hd__clkbuf_4 T11Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5303));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R0_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5339));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R1_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R2_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R2_INV_1 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5375));
  sky130_fd_sc_hd__clkbuf_4 T11Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B444));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R0_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y4__R1_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B30));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R1_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R2_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R2_INV_1 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B516));
  sky130_fd_sc_hd__clkbuf_4 T11Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5411));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R0_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5447));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R1_INV_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R2_INV_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R2_INV_1 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5483));
  sky130_fd_sc_hd__clkbuf_4 T11Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5519));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R0_INV_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5555));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R1_INV_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R2_INV_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R2_INV_1 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5591));
  sky130_fd_sc_hd__clkbuf_4 T11Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5627));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R0_INV_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5663));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R1_INV_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R2_INV_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R2_INV_1 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5699));
  sky130_fd_sc_hd__clkbuf_4 T11Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5735));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R0_INV_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5771));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R1_INV_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R2_INV_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R2_INV_1 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5807));
  sky130_fd_sc_hd__clkbuf_4 T11Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5843));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R0_INV_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5879));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R1_INV_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R2_INV_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R2_INV_1 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5915));
  sky130_fd_sc_hd__clkbuf_4 T11Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5951));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R0_INV_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5987));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R1_INV_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R2_INV_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R2_INV_1 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6023));
  sky130_fd_sc_hd__clkbuf_4 T11Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6059));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R0_INV_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6095));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R1_INV_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R2_INV_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R2_INV_1 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6131));
  sky130_fd_sc_hd__clkbuf_4 T11Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6167));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R0_INV_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6203));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R1_INV_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R2_INV_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R2_INV_1 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6239));
  sky130_fd_sc_hd__clkbuf_4 T11Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6275));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R0_INV_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6311));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R1_INV_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R2_INV_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R2_INV_1 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6347));
  sky130_fd_sc_hd__clkbuf_4 T11Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6383));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R0_INV_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6419));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R1_INV_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R2_INV_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R2_INV_1 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6455));
  sky130_fd_sc_hd__clkbuf_4 T11Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B552));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R0_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B588));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R1_INV_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R2_INV_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R2_INV_1 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y5__R3_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B39));
  sky130_fd_sc_hd__clkbuf_4 T11Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6491));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R0_INV_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6527));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R1_INV_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R2_INV_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R2_INV_1 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6563));
  sky130_fd_sc_hd__clkbuf_4 T11Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6599));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R0_INV_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6635));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R1_INV_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R2_INV_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R2_INV_1 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6671));
  sky130_fd_sc_hd__clkbuf_4 T11Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6707));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R0_INV_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6743));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R1_INV_0 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R2_INV_0 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R2_INV_1 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6779));
  sky130_fd_sc_hd__clkbuf_4 T11Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6815));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R0_INV_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6851));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R1_INV_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R2_INV_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R2_INV_1 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6887));
  sky130_fd_sc_hd__clkbuf_4 T11Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6923));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R0_INV_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6959));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R1_INV_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R2_INV_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R2_INV_1 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6995));
  sky130_fd_sc_hd__clkbuf_4 T11Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7031));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R0_INV_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7067));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R1_INV_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R2_INV_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R2_INV_1 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7103));
  sky130_fd_sc_hd__clkbuf_4 T11Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7139));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R0_INV_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7175));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R1_INV_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R2_INV_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R2_INV_1 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7211));
  sky130_fd_sc_hd__clkbuf_4 T11Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7247));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R0_INV_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7283));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R1_INV_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R2_INV_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R2_INV_1 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7319));
  sky130_fd_sc_hd__clkbuf_4 T11Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7355));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R0_INV_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7391));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R1_INV_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R2_INV_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R2_INV_1 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7427));
  sky130_fd_sc_hd__clkbuf_4 T11Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7463));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R0_INV_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7499));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R1_INV_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R2_INV_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R2_INV_1 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7535));
  sky130_fd_sc_hd__clkbuf_4 T11Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B660));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R0_INV_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B696));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R1_INV_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R2_INV_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R2_INV_1 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B732));
  sky130_fd_sc_hd__clkbuf_4 T11Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7571));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R0_INV_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7607));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R1_INV_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R2_INV_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R2_INV_1 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7643));
  sky130_fd_sc_hd__clkbuf_4 T11Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7679));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R0_INV_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7715));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R1_INV_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R2_INV_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R2_INV_1 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7751));
  sky130_fd_sc_hd__clkbuf_4 T11Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7787));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R0_INV_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7823));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R1_INV_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R2_INV_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R2_INV_1 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7859));
  sky130_fd_sc_hd__clkbuf_4 T11Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7895));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R0_INV_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7931));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R1_INV_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R2_INV_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R2_INV_1 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7967));
  sky130_fd_sc_hd__clkbuf_4 T11Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8003));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R0_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8039));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R1_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R2_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R2_INV_1 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8075));
  sky130_fd_sc_hd__clkbuf_4 T11Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8111));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R0_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8147));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R1_INV_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R2_INV_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R2_INV_1 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8183));
  sky130_fd_sc_hd__clkbuf_4 T11Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8219));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R0_INV_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8255));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R1_INV_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R2_INV_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R2_INV_1 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8291));
  sky130_fd_sc_hd__clkbuf_4 T11Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8327));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R0_INV_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8363));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R1_INV_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R2_INV_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R2_INV_1 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8399));
  sky130_fd_sc_hd__clkbuf_4 T11Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8435));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R0_INV_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8471));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R1_INV_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R2_INV_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R2_INV_1 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8507));
  sky130_fd_sc_hd__clkbuf_4 T11Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8543));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R0_INV_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8579));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R1_INV_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R2_INV_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R2_INV_1 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8615));
  sky130_fd_sc_hd__clkbuf_4 T11Y7__R0_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B3));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R0_INV_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B804));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R1_INV_0 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R2_INV_0 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R2_INV_1 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B840));
  sky130_fd_sc_hd__clkbuf_4 T11Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8651));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R0_INV_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8687));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R1_INV_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R2_INV_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R2_INV_1 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8723));
  sky130_fd_sc_hd__clkbuf_4 T11Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8759));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R0_INV_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8795));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R1_INV_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R2_INV_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R2_INV_1 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8831));
  sky130_fd_sc_hd__clkbuf_4 T11Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8867));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R0_INV_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8903));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R1_INV_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R2_INV_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R2_INV_1 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8939));
  sky130_fd_sc_hd__clkbuf_4 T11Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8975));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R0_INV_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9011));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R1_INV_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R2_INV_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R2_INV_1 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9047));
  sky130_fd_sc_hd__clkbuf_4 T11Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9083));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R0_INV_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9119));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R1_INV_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R2_INV_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R2_INV_1 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9155));
  sky130_fd_sc_hd__clkbuf_4 T11Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9191));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R0_INV_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9227));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R1_INV_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R2_INV_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R2_INV_1 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9263));
  sky130_fd_sc_hd__clkbuf_4 T11Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9299));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R0_INV_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9335));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R1_INV_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R2_INV_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R2_INV_1 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9371));
  sky130_fd_sc_hd__clkbuf_4 T11Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9407));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R0_INV_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9443));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R1_INV_0 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R2_INV_0 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R2_INV_1 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9479));
  sky130_fd_sc_hd__clkbuf_4 T11Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9515));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R0_INV_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9551));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R1_INV_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R2_INV_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R2_INV_1 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9587));
  sky130_fd_sc_hd__clkbuf_4 T11Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9623));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R0_INV_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9659));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R1_INV_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R2_INV_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R2_INV_1 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9695));
  sky130_fd_sc_hd__clkbuf_4 T11Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B876));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R0_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y8__R1_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B57));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R1_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R2_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R2_INV_1 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B948));
  sky130_fd_sc_hd__clkbuf_4 T11Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B984));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R0_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1020));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R1_INV_0 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R2_INV_0 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R2_INV_1 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y9__R3_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B66));
  sky130_fd_sc_hd__clkbuf_4 T12Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B22));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R0_INV_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B57));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R1_INV_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R2_INV_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R2_INV_1 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B92));
  sky130_fd_sc_hd__clkbuf_4 T12Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1093));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R0_INV_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1129));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R1_INV_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R2_INV_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R2_INV_1 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1165));
  sky130_fd_sc_hd__clkbuf_4 T12Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1201));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R0_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1237));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R1_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R2_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R2_INV_1 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1273));
  sky130_fd_sc_hd__clkbuf_4 T12Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1309));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R0_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1345));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R1_INV_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R2_INV_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R2_INV_1 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1381));
  sky130_fd_sc_hd__clkbuf_4 T12Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1417));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R0_INV_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1453));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R1_INV_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R2_INV_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R2_INV_1 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1489));
  sky130_fd_sc_hd__clkbuf_4 T12Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1525));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R0_INV_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1560));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R1_INV_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R2_INV_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R2_INV_1 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1596));
  sky130_fd_sc_hd__clkbuf_4 T12Y15__R0_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B102));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R0_INV_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1668));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R1_INV_0 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R2_INV_0 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R2_INV_1 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1704));
  sky130_fd_sc_hd__clkbuf_4 T12Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1740));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R0_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y16__R1_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B111));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R1_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R2_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R2_INV_1 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1812));
  sky130_fd_sc_hd__clkbuf_4 T12Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1848));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R0_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1884));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R1_INV_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R2_INV_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R2_INV_1 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y17__R3_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B120));
  sky130_fd_sc_hd__clkbuf_4 T12Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1956));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R0_INV_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1992));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R1_INV_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R2_INV_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R2_INV_1 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2028));
  sky130_fd_sc_hd__clkbuf_4 T12Y19__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B129));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R0_INV_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2100));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R1_INV_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R2_INV_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R2_INV_1 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2136));
  sky130_fd_sc_hd__clkbuf_4 T12Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B127));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R0_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B162));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R1_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R2_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R2_INV_1 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B197));
  sky130_fd_sc_hd__clkbuf_4 T12Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2172));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R0_INV_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y20__R1_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B138));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R1_INV_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R2_INV_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R2_INV_1 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2244));
  sky130_fd_sc_hd__clkbuf_4 T12Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2280));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R0_INV_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2316));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R1_INV_0 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R2_INV_0 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R2_INV_1 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y21__R3_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B147));
  sky130_fd_sc_hd__clkbuf_4 T12Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2388));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R0_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2424));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R1_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R2_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R2_INV_1 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2460));
  sky130_fd_sc_hd__clkbuf_4 T12Y23__R0_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B156));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R0_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2532));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R1_INV_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R2_INV_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R2_INV_1 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2568));
  sky130_fd_sc_hd__clkbuf_4 T12Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2604));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R0_INV_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y24__R1_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B165));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R1_INV_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R2_INV_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R2_INV_1 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2676));
  sky130_fd_sc_hd__clkbuf_4 T12Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2712));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R0_INV_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2748));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R1_INV_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R2_INV_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R2_INV_1 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y25__R3_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B174));
  sky130_fd_sc_hd__clkbuf_4 T12Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2820));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R0_INV_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2856));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R1_INV_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R2_INV_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R2_INV_1 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2892));
  sky130_fd_sc_hd__clkbuf_4 T12Y27__R0_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B183));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R0_INV_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2964));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R1_INV_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R2_INV_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R2_INV_1 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3000));
  sky130_fd_sc_hd__clkbuf_4 T12Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3036));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R0_INV_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y28__R1_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B12));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R1_INV_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R2_INV_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R2_INV_1 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3108));
  sky130_fd_sc_hd__clkbuf_4 T12Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3144));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R0_INV_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3180));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R1_INV_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R2_INV_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R2_INV_1 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y29__R3_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B201));
  sky130_fd_sc_hd__clkbuf_4 T12Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B232));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R0_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B267));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R1_INV_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R2_INV_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R2_INV_1 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B303));
  sky130_fd_sc_hd__clkbuf_4 T12Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3252));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R0_INV_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3288));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R1_INV_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R2_INV_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R2_INV_1 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3324));
  sky130_fd_sc_hd__clkbuf_4 T12Y31__R0_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B210));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R0_INV_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3396));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R1_INV_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R2_INV_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R2_INV_1 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3432));
  sky130_fd_sc_hd__clkbuf_4 T12Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3468));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R0_INV_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y32__R1_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B219));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R1_INV_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R2_INV_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R2_INV_1 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3540));
  sky130_fd_sc_hd__clkbuf_4 T12Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3576));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R0_INV_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3612));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R1_INV_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R2_INV_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R2_INV_1 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y33__R3_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B228));
  sky130_fd_sc_hd__clkbuf_4 T12Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3684));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R0_INV_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3720));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R1_INV_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R2_INV_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R2_INV_1 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3756));
  sky130_fd_sc_hd__clkbuf_4 T12Y35__R0_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B237));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R0_INV_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3828));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R1_INV_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R2_INV_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R2_INV_1 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3864));
  sky130_fd_sc_hd__clkbuf_4 T12Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3900));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R0_INV_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y36__R1_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B246));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R1_INV_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R2_INV_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R2_INV_1 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3972));
  sky130_fd_sc_hd__clkbuf_4 T12Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4008));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R0_INV_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4044));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R1_INV_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R2_INV_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R2_INV_1 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y37__R3_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B255));
  sky130_fd_sc_hd__clkbuf_4 T12Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4116));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R0_INV_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4152));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R1_INV_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R2_INV_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R2_INV_1 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4188));
  sky130_fd_sc_hd__clkbuf_4 T12Y39__R0_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B264));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R0_INV_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4260));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R1_INV_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R2_INV_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R2_INV_1 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4296));
  sky130_fd_sc_hd__clkbuf_4 T12Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B338));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R0_INV_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B373));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R1_INV_0 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R2_INV_0 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R2_INV_1 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B409));
  sky130_fd_sc_hd__clkbuf_4 T12Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4332));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R0_INV_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y40__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B273));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R1_INV_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R2_INV_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R2_INV_1 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4404));
  sky130_fd_sc_hd__clkbuf_4 T12Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4440));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R0_INV_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4476));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R1_INV_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R2_INV_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R2_INV_1 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y41__R3_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B282));
  sky130_fd_sc_hd__clkbuf_4 T12Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4548));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R0_INV_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4584));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R1_INV_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R2_INV_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R2_INV_1 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4620));
  sky130_fd_sc_hd__clkbuf_4 T12Y43__R0_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B291));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R0_INV_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4692));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R1_INV_0 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R2_INV_0 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R2_INV_1 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4728));
  sky130_fd_sc_hd__clkbuf_4 T12Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4764));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R0_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y44__R1_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B300));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R1_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R2_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R2_INV_1 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4836));
  sky130_fd_sc_hd__clkbuf_4 T12Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4872));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R0_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4908));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R1_INV_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R2_INV_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R2_INV_1 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y45__R3_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B309));
  sky130_fd_sc_hd__clkbuf_4 T12Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4980));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R0_INV_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5016));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R1_INV_0 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R2_INV_0 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R2_INV_1 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5052));
  sky130_fd_sc_hd__clkbuf_4 T12Y47__R0_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B318));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R0_INV_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5124));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R1_INV_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R2_INV_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R2_INV_1 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5160));
  sky130_fd_sc_hd__clkbuf_4 T12Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5196));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R0_INV_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y48__R1_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B327));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R1_INV_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R2_INV_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R2_INV_1 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5268));
  sky130_fd_sc_hd__clkbuf_4 T12Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5304));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R0_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5340));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R1_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R2_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R2_INV_1 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y49__R3_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B21));
  sky130_fd_sc_hd__clkbuf_4 T12Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B445));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R0_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B481));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R1_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R2_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R2_INV_1 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B517));
  sky130_fd_sc_hd__clkbuf_4 T12Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5412));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R0_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5448));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R1_INV_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R2_INV_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R2_INV_1 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5484));
  sky130_fd_sc_hd__clkbuf_4 T12Y51__R0_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B345));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R0_INV_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5556));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R1_INV_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R2_INV_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R2_INV_1 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5592));
  sky130_fd_sc_hd__clkbuf_4 T12Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5628));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R0_INV_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y52__R1_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B354));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R1_INV_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R2_INV_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R2_INV_1 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5700));
  sky130_fd_sc_hd__clkbuf_4 T12Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5736));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R0_INV_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5772));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R1_INV_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R2_INV_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R2_INV_1 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y53__R3_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B363));
  sky130_fd_sc_hd__clkbuf_4 T12Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5844));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R0_INV_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5880));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R1_INV_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R2_INV_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R2_INV_1 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5916));
  sky130_fd_sc_hd__clkbuf_4 T12Y55__R0_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B372));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R0_INV_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5988));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R1_INV_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R2_INV_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R2_INV_1 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6024));
  sky130_fd_sc_hd__clkbuf_4 T12Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6060));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R0_INV_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y56__R1_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B381));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R1_INV_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R2_INV_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R2_INV_1 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6132));
  sky130_fd_sc_hd__clkbuf_4 T12Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6168));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R0_INV_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6204));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R1_INV_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R2_INV_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R2_INV_1 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y57__R3_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B390));
  sky130_fd_sc_hd__clkbuf_4 T12Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6276));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R0_INV_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6312));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R1_INV_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R2_INV_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R2_INV_1 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6348));
  sky130_fd_sc_hd__clkbuf_4 T12Y59__R0_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B399));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R0_INV_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6420));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R1_INV_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R2_INV_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R2_INV_1 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6456));
  sky130_fd_sc_hd__clkbuf_4 T12Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B553));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R0_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B589));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R1_INV_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R2_INV_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R2_INV_1 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B625));
  sky130_fd_sc_hd__clkbuf_4 T12Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6492));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R0_INV_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y60__R1_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B408));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R1_INV_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R2_INV_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R2_INV_1 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6564));
  sky130_fd_sc_hd__clkbuf_4 T12Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6600));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R0_INV_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6636));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R1_INV_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R2_INV_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R2_INV_1 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y61__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B417));
  sky130_fd_sc_hd__clkbuf_4 T12Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6708));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R0_INV_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6744));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R1_INV_0 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R2_INV_0 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R2_INV_1 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6780));
  sky130_fd_sc_hd__clkbuf_4 T12Y63__R0_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B426));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R0_INV_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6852));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R1_INV_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R2_INV_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R2_INV_1 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6888));
  sky130_fd_sc_hd__clkbuf_4 T12Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6924));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R0_INV_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y64__R1_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B435));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R1_INV_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R2_INV_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R2_INV_1 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6996));
  sky130_fd_sc_hd__clkbuf_4 T12Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7032));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R0_INV_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7068));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R1_INV_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R2_INV_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R2_INV_1 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y65__R3_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B444));
  sky130_fd_sc_hd__clkbuf_4 T12Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7140));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R0_INV_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7176));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R1_INV_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R2_INV_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R2_INV_1 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7212));
  sky130_fd_sc_hd__clkbuf_4 T12Y67__R0_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B453));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R0_INV_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7284));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R1_INV_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R2_INV_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R2_INV_1 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7320));
  sky130_fd_sc_hd__clkbuf_4 T12Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7356));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R0_INV_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y68__R1_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B462));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R1_INV_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R2_INV_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R2_INV_1 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7428));
  sky130_fd_sc_hd__clkbuf_4 T12Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7464));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R0_INV_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7500));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R1_INV_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R2_INV_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R2_INV_1 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y69__R3_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B471));
  sky130_fd_sc_hd__clkbuf_4 T12Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B661));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R0_INV_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B697));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R1_INV_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R2_INV_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R2_INV_1 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B733));
  sky130_fd_sc_hd__clkbuf_4 T12Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7572));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R0_INV_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7608));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R1_INV_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R2_INV_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R2_INV_1 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7644));
  sky130_fd_sc_hd__clkbuf_4 T12Y71__R0_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B30));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R0_INV_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7716));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R1_INV_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R2_INV_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R2_INV_1 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7752));
  sky130_fd_sc_hd__clkbuf_4 T12Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7788));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R0_INV_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y72__R1_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B489));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R1_INV_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R2_INV_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R2_INV_1 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7860));
  sky130_fd_sc_hd__clkbuf_4 T12Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7896));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R0_INV_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7932));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R1_INV_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R2_INV_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R2_INV_1 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y73__R3_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B498));
  sky130_fd_sc_hd__clkbuf_4 T12Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8004));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R0_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8040));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R1_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R2_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R2_INV_1 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8076));
  sky130_fd_sc_hd__clkbuf_4 T12Y75__R0_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B507));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R0_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8148));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R1_INV_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R2_INV_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R2_INV_1 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8184));
  sky130_fd_sc_hd__clkbuf_4 T12Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8220));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R0_INV_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y76__R1_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B516));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R1_INV_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R2_INV_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R2_INV_1 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8292));
  sky130_fd_sc_hd__clkbuf_4 T12Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8328));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R0_INV_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8364));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R1_INV_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R2_INV_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R2_INV_1 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y77__R3_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B525));
  sky130_fd_sc_hd__clkbuf_4 T12Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8436));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R0_INV_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8472));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R1_INV_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R2_INV_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R2_INV_1 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8508));
  sky130_fd_sc_hd__clkbuf_4 T12Y79__R0_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B534));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R0_INV_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8580));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R1_INV_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R2_INV_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R2_INV_1 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8616));
  sky130_fd_sc_hd__clkbuf_4 T12Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B769));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R0_INV_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B805));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R1_INV_0 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R2_INV_0 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R2_INV_1 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B841));
  sky130_fd_sc_hd__clkbuf_4 T12Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8652));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R0_INV_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y80__R1_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B543));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R1_INV_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R2_INV_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R2_INV_1 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8724));
  sky130_fd_sc_hd__clkbuf_4 T12Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8760));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R0_INV_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8796));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R1_INV_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R2_INV_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R2_INV_1 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y81__R3_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B552));
  sky130_fd_sc_hd__clkbuf_4 T12Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8868));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R0_INV_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8904));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R1_INV_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R2_INV_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R2_INV_1 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8940));
  sky130_fd_sc_hd__clkbuf_4 T12Y83__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B561));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R0_INV_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9012));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R1_INV_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R2_INV_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R2_INV_1 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9048));
  sky130_fd_sc_hd__clkbuf_4 T12Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9084));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R0_INV_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y84__R1_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B570));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R1_INV_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R2_INV_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R2_INV_1 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9156));
  sky130_fd_sc_hd__clkbuf_4 T12Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9192));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R0_INV_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9228));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R1_INV_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R2_INV_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R2_INV_1 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y85__R3_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B579));
  sky130_fd_sc_hd__clkbuf_4 T12Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9300));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R0_INV_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9336));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R1_INV_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R2_INV_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R2_INV_1 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9372));
  sky130_fd_sc_hd__clkbuf_4 T12Y87__R0_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B588));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R0_INV_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9444));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R1_INV_0 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R2_INV_0 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R2_INV_1 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9480));
  sky130_fd_sc_hd__clkbuf_4 T12Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9516));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R0_INV_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y88__R1_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B597));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R1_INV_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R2_INV_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R2_INV_1 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9588));
  sky130_fd_sc_hd__clkbuf_4 T12Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9624));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R0_INV_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9660));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R1_INV_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R2_INV_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R2_INV_1 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y89__R3_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B606));
  sky130_fd_sc_hd__clkbuf_4 T12Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B877));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R0_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B913));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R1_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R2_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R2_INV_1 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B949));
  sky130_fd_sc_hd__clkbuf_4 T12Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B985));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R0_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1021));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R1_INV_0 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R2_INV_0 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R2_INV_1 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1057));
  sky130_fd_sc_hd__clkbuf_4 T13Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B23));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R0_INV_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B58));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R1_INV_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R2_INV_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R2_INV_1 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B93));
  sky130_fd_sc_hd__clkbuf_4 T13Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1094));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R0_INV_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1130));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R1_INV_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R2_INV_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R2_INV_1 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1166));
  sky130_fd_sc_hd__clkbuf_4 T13Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1202));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R0_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1238));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R1_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R2_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R2_INV_1 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1274));
  sky130_fd_sc_hd__clkbuf_4 T13Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1310));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R0_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1346));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R1_INV_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R2_INV_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R2_INV_1 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1382));
  sky130_fd_sc_hd__clkbuf_4 T13Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1418));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R0_INV_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1454));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R1_INV_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R2_INV_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R2_INV_1 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1490));
  sky130_fd_sc_hd__clkbuf_4 T13Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1526));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R0_INV_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1561));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R1_INV_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R2_INV_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R2_INV_1 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1597));
  sky130_fd_sc_hd__clkbuf_4 T13Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1633));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R0_INV_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1669));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R1_INV_0 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R2_INV_0 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R2_INV_1 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1705));
  sky130_fd_sc_hd__clkbuf_4 T13Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1741));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R0_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1777));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R1_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R2_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R2_INV_1 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1813));
  sky130_fd_sc_hd__clkbuf_4 T13Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1849));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R0_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1885));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R1_INV_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R2_INV_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R2_INV_1 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1921));
  sky130_fd_sc_hd__clkbuf_4 T13Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1957));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R0_INV_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1993));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R1_INV_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R2_INV_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R2_INV_1 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2029));
  sky130_fd_sc_hd__clkbuf_4 T13Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2065));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R0_INV_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2101));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R1_INV_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R2_INV_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R2_INV_1 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2137));
  sky130_fd_sc_hd__clkbuf_4 T13Y1__R0_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B8));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R0_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B163));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R1_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R2_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R2_INV_1 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B198));
  sky130_fd_sc_hd__clkbuf_4 T13Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2173));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R0_INV_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2209));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R1_INV_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R2_INV_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R2_INV_1 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2245));
  sky130_fd_sc_hd__clkbuf_4 T13Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2281));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R0_INV_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2317));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R1_INV_0 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R2_INV_0 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R2_INV_1 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2353));
  sky130_fd_sc_hd__clkbuf_4 T13Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2389));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R0_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2425));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R1_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R2_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R2_INV_1 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2461));
  sky130_fd_sc_hd__clkbuf_4 T13Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2497));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R0_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2533));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R1_INV_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R2_INV_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R2_INV_1 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2569));
  sky130_fd_sc_hd__clkbuf_4 T13Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2605));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R0_INV_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2641));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R1_INV_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R2_INV_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R2_INV_1 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2677));
  sky130_fd_sc_hd__clkbuf_4 T13Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2713));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R0_INV_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2749));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R1_INV_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R2_INV_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R2_INV_1 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2785));
  sky130_fd_sc_hd__clkbuf_4 T13Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2821));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R0_INV_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2857));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R1_INV_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R2_INV_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R2_INV_1 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2893));
  sky130_fd_sc_hd__clkbuf_4 T13Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2929));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R0_INV_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2965));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R1_INV_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R2_INV_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R2_INV_1 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3001));
  sky130_fd_sc_hd__clkbuf_4 T13Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3037));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R0_INV_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3073));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R1_INV_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R2_INV_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R2_INV_1 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3109));
  sky130_fd_sc_hd__clkbuf_4 T13Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3145));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R0_INV_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3181));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R1_INV_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R2_INV_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R2_INV_1 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3217));
  sky130_fd_sc_hd__clkbuf_4 T13Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B233));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R0_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B268));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R1_INV_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R2_INV_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R2_INV_1 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y2__R3_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B19));
  sky130_fd_sc_hd__clkbuf_4 T13Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3253));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R0_INV_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3289));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R1_INV_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R2_INV_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R2_INV_1 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3325));
  sky130_fd_sc_hd__clkbuf_4 T13Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3361));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R0_INV_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3397));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R1_INV_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R2_INV_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R2_INV_1 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3433));
  sky130_fd_sc_hd__clkbuf_4 T13Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3469));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R0_INV_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3505));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R1_INV_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R2_INV_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R2_INV_1 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3541));
  sky130_fd_sc_hd__clkbuf_4 T13Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3577));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R0_INV_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3613));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R1_INV_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R2_INV_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R2_INV_1 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3649));
  sky130_fd_sc_hd__clkbuf_4 T13Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3685));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R0_INV_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3721));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R1_INV_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R2_INV_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R2_INV_1 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3757));
  sky130_fd_sc_hd__clkbuf_4 T13Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3793));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R0_INV_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3829));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R1_INV_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R2_INV_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R2_INV_1 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3865));
  sky130_fd_sc_hd__clkbuf_4 T13Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3901));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R0_INV_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3937));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R1_INV_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R2_INV_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R2_INV_1 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3973));
  sky130_fd_sc_hd__clkbuf_4 T13Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4009));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R0_INV_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4045));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R1_INV_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R2_INV_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R2_INV_1 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4081));
  sky130_fd_sc_hd__clkbuf_4 T13Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4117));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R0_INV_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4153));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R1_INV_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R2_INV_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R2_INV_1 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4189));
  sky130_fd_sc_hd__clkbuf_4 T13Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4225));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R0_INV_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4261));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R1_INV_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R2_INV_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R2_INV_1 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4297));
  sky130_fd_sc_hd__clkbuf_4 T13Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B339));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R0_INV_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B374));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R1_INV_0 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R2_INV_0 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R2_INV_1 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B410));
  sky130_fd_sc_hd__clkbuf_4 T13Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4333));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R0_INV_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4369));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R1_INV_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R2_INV_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R2_INV_1 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4405));
  sky130_fd_sc_hd__clkbuf_4 T13Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4441));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R0_INV_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4477));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R1_INV_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R2_INV_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R2_INV_1 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4513));
  sky130_fd_sc_hd__clkbuf_4 T13Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4549));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R0_INV_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4585));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R1_INV_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R2_INV_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R2_INV_1 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4621));
  sky130_fd_sc_hd__clkbuf_4 T13Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4657));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R0_INV_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4693));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R1_INV_0 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R2_INV_0 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R2_INV_1 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4729));
  sky130_fd_sc_hd__clkbuf_4 T13Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4765));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R0_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4801));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R1_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R2_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R2_INV_1 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4837));
  sky130_fd_sc_hd__clkbuf_4 T13Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4873));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R0_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4909));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R1_INV_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R2_INV_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R2_INV_1 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4945));
  sky130_fd_sc_hd__clkbuf_4 T13Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4981));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R0_INV_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5017));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R1_INV_0 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R2_INV_0 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R2_INV_1 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5053));
  sky130_fd_sc_hd__clkbuf_4 T13Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5089));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R0_INV_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5125));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R1_INV_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R2_INV_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R2_INV_1 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5161));
  sky130_fd_sc_hd__clkbuf_4 T13Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5197));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R0_INV_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5233));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R1_INV_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R2_INV_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R2_INV_1 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5269));
  sky130_fd_sc_hd__clkbuf_4 T13Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5305));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R0_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5341));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R1_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R2_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R2_INV_1 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5377));
  sky130_fd_sc_hd__clkbuf_4 T13Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B446));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R0_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B482));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R1_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R2_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R2_INV_1 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B518));
  sky130_fd_sc_hd__clkbuf_4 T13Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5413));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R0_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5449));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R1_INV_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R2_INV_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R2_INV_1 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5485));
  sky130_fd_sc_hd__clkbuf_4 T13Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5521));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R0_INV_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5557));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R1_INV_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R2_INV_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R2_INV_1 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5593));
  sky130_fd_sc_hd__clkbuf_4 T13Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5629));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R0_INV_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5665));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R1_INV_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R2_INV_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R2_INV_1 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5701));
  sky130_fd_sc_hd__clkbuf_4 T13Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5737));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R0_INV_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5773));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R1_INV_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R2_INV_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R2_INV_1 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5809));
  sky130_fd_sc_hd__clkbuf_4 T13Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5845));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R0_INV_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5881));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R1_INV_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R2_INV_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R2_INV_1 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5917));
  sky130_fd_sc_hd__clkbuf_4 T13Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5953));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R0_INV_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5989));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R1_INV_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R2_INV_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R2_INV_1 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6025));
  sky130_fd_sc_hd__clkbuf_4 T13Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6061));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R0_INV_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6097));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R1_INV_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R2_INV_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R2_INV_1 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6133));
  sky130_fd_sc_hd__clkbuf_4 T13Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6169));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R0_INV_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6205));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R1_INV_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R2_INV_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R2_INV_1 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6241));
  sky130_fd_sc_hd__clkbuf_4 T13Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6277));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R0_INV_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6313));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R1_INV_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R2_INV_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R2_INV_1 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6349));
  sky130_fd_sc_hd__clkbuf_4 T13Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6385));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R0_INV_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6421));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R1_INV_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R2_INV_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R2_INV_1 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6457));
  sky130_fd_sc_hd__clkbuf_4 T13Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B554));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R0_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B590));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R1_INV_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R2_INV_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R2_INV_1 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B626));
  sky130_fd_sc_hd__clkbuf_4 T13Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6493));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R0_INV_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6529));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R1_INV_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R2_INV_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R2_INV_1 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6565));
  sky130_fd_sc_hd__clkbuf_4 T13Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6601));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R0_INV_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6637));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R1_INV_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R2_INV_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R2_INV_1 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6673));
  sky130_fd_sc_hd__clkbuf_4 T13Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6709));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R0_INV_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6745));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R1_INV_0 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R2_INV_0 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R2_INV_1 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6781));
  sky130_fd_sc_hd__clkbuf_4 T13Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6817));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R0_INV_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6853));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R1_INV_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R2_INV_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R2_INV_1 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6889));
  sky130_fd_sc_hd__clkbuf_4 T13Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6925));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R0_INV_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6961));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R1_INV_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R2_INV_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R2_INV_1 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6997));
  sky130_fd_sc_hd__clkbuf_4 T13Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7033));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R0_INV_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7069));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R1_INV_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R2_INV_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R2_INV_1 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7105));
  sky130_fd_sc_hd__clkbuf_4 T13Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7141));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R0_INV_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7177));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R1_INV_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R2_INV_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R2_INV_1 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7213));
  sky130_fd_sc_hd__clkbuf_4 T13Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7249));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R0_INV_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7285));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R1_INV_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R2_INV_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R2_INV_1 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7321));
  sky130_fd_sc_hd__clkbuf_4 T13Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7357));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R0_INV_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7393));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R1_INV_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R2_INV_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R2_INV_1 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7429));
  sky130_fd_sc_hd__clkbuf_4 T13Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7465));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R0_INV_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7501));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R1_INV_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R2_INV_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R2_INV_1 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7537));
  sky130_fd_sc_hd__clkbuf_4 T13Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B662));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R0_INV_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B698));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R1_INV_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R2_INV_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R2_INV_1 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B734));
  sky130_fd_sc_hd__clkbuf_4 T13Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7573));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R0_INV_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7609));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R1_INV_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R2_INV_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R2_INV_1 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7645));
  sky130_fd_sc_hd__clkbuf_4 T13Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7681));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R0_INV_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7717));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R1_INV_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R2_INV_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R2_INV_1 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7753));
  sky130_fd_sc_hd__clkbuf_4 T13Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7789));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R0_INV_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7825));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R1_INV_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R2_INV_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R2_INV_1 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7861));
  sky130_fd_sc_hd__clkbuf_4 T13Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7897));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R0_INV_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7933));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R1_INV_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R2_INV_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R2_INV_1 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7969));
  sky130_fd_sc_hd__clkbuf_4 T13Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8005));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R0_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8041));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R1_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R2_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R2_INV_1 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8077));
  sky130_fd_sc_hd__clkbuf_4 T13Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8113));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R0_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8149));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R1_INV_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R2_INV_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R2_INV_1 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8185));
  sky130_fd_sc_hd__clkbuf_4 T13Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8221));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R0_INV_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8257));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R1_INV_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R2_INV_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R2_INV_1 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8293));
  sky130_fd_sc_hd__clkbuf_4 T13Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8329));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R0_INV_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8365));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R1_INV_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R2_INV_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R2_INV_1 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8401));
  sky130_fd_sc_hd__clkbuf_4 T13Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8437));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R0_INV_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8473));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R1_INV_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R2_INV_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R2_INV_1 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8509));
  sky130_fd_sc_hd__clkbuf_4 T13Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8545));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R0_INV_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8581));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R1_INV_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R2_INV_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R2_INV_1 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8617));
  sky130_fd_sc_hd__clkbuf_4 T13Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B770));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R0_INV_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B806));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R1_INV_0 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R2_INV_0 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R2_INV_1 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B842));
  sky130_fd_sc_hd__clkbuf_4 T13Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8653));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R0_INV_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8689));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R1_INV_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R2_INV_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R2_INV_1 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8725));
  sky130_fd_sc_hd__clkbuf_4 T13Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8761));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R0_INV_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8797));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R1_INV_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R2_INV_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R2_INV_1 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8833));
  sky130_fd_sc_hd__clkbuf_4 T13Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8869));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R0_INV_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8905));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R1_INV_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R2_INV_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R2_INV_1 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8941));
  sky130_fd_sc_hd__clkbuf_4 T13Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8977));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R0_INV_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9013));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R1_INV_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R2_INV_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R2_INV_1 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9049));
  sky130_fd_sc_hd__clkbuf_4 T13Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9085));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R0_INV_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9121));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R1_INV_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R2_INV_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R2_INV_1 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9157));
  sky130_fd_sc_hd__clkbuf_4 T13Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9193));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R0_INV_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9229));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R1_INV_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R2_INV_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R2_INV_1 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9265));
  sky130_fd_sc_hd__clkbuf_4 T13Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9301));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R0_INV_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9337));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R1_INV_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R2_INV_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R2_INV_1 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9373));
  sky130_fd_sc_hd__clkbuf_4 T13Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9409));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R0_INV_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9445));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R1_INV_0 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R2_INV_0 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R2_INV_1 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9481));
  sky130_fd_sc_hd__clkbuf_4 T13Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9517));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R0_INV_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9553));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R1_INV_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R2_INV_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R2_INV_1 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9589));
  sky130_fd_sc_hd__clkbuf_4 T13Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9625));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R0_INV_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9661));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R1_INV_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R2_INV_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R2_INV_1 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9697));
  sky130_fd_sc_hd__clkbuf_4 T13Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B878));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R0_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B914));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R1_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R2_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R2_INV_1 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B950));
  sky130_fd_sc_hd__clkbuf_4 T13Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B986));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R0_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1022));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R1_INV_0 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R2_INV_0 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R2_INV_1 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1058));
  sky130_fd_sc_hd__clkbuf_4 T14Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B24));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R0_INV_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B59));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R1_INV_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R2_INV_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R2_INV_1 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B94));
  sky130_fd_sc_hd__clkbuf_4 T14Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1095));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R0_INV_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1131));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R1_INV_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R2_INV_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R2_INV_1 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1167));
  sky130_fd_sc_hd__clkbuf_4 T14Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1203));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R0_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1239));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R1_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R2_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R2_INV_1 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1275));
  sky130_fd_sc_hd__clkbuf_4 T14Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1311));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R0_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1347));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R1_INV_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R2_INV_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R2_INV_1 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1383));
  sky130_fd_sc_hd__clkbuf_4 T14Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1419));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R0_INV_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1455));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R1_INV_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R2_INV_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R2_INV_1 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1491));
  sky130_fd_sc_hd__clkbuf_4 T14Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1527));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R0_INV_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1562));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R1_INV_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R2_INV_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R2_INV_1 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1598));
  sky130_fd_sc_hd__clkbuf_4 T14Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1634));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R0_INV_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1670));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R1_INV_0 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R2_INV_0 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R2_INV_1 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1706));
  sky130_fd_sc_hd__clkbuf_4 T14Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1742));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R0_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1778));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R1_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R2_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R2_INV_1 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1814));
  sky130_fd_sc_hd__clkbuf_4 T14Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1850));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R0_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1886));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R1_INV_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R2_INV_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R2_INV_1 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1922));
  sky130_fd_sc_hd__clkbuf_4 T14Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1958));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R0_INV_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1994));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R1_INV_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R2_INV_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R2_INV_1 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2030));
  sky130_fd_sc_hd__clkbuf_4 T14Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2066));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R0_INV_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2102));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R1_INV_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R2_INV_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R2_INV_1 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2138));
  sky130_fd_sc_hd__clkbuf_4 T14Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B129));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R0_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B164));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R1_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R2_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R2_INV_1 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B199));
  sky130_fd_sc_hd__clkbuf_4 T14Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2174));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R0_INV_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2210));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R1_INV_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R2_INV_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R2_INV_1 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2246));
  sky130_fd_sc_hd__clkbuf_4 T14Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2282));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R0_INV_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2318));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R1_INV_0 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R2_INV_0 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R2_INV_1 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2354));
  sky130_fd_sc_hd__clkbuf_4 T14Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2390));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R0_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2426));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R1_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R2_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R2_INV_1 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2462));
  sky130_fd_sc_hd__clkbuf_4 T14Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2498));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R0_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2534));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R1_INV_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R2_INV_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R2_INV_1 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2570));
  sky130_fd_sc_hd__clkbuf_4 T14Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2606));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R0_INV_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2642));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R1_INV_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R2_INV_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R2_INV_1 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2678));
  sky130_fd_sc_hd__clkbuf_4 T14Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2714));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R0_INV_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2750));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R1_INV_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R2_INV_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R2_INV_1 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2786));
  sky130_fd_sc_hd__clkbuf_4 T14Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2822));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R0_INV_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2858));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R1_INV_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R2_INV_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R2_INV_1 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2894));
  sky130_fd_sc_hd__clkbuf_4 T14Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2930));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R0_INV_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2966));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R1_INV_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R2_INV_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R2_INV_1 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3002));
  sky130_fd_sc_hd__clkbuf_4 T14Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3038));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R0_INV_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3074));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R1_INV_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R2_INV_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R2_INV_1 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3110));
  sky130_fd_sc_hd__clkbuf_4 T14Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3146));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R0_INV_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3182));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R1_INV_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R2_INV_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R2_INV_1 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3218));
  sky130_fd_sc_hd__clkbuf_4 T14Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B234));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R0_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B269));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R1_INV_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R2_INV_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R2_INV_1 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B305));
  sky130_fd_sc_hd__clkbuf_4 T14Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3254));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R0_INV_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3290));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R1_INV_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R2_INV_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R2_INV_1 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3326));
  sky130_fd_sc_hd__clkbuf_4 T14Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3362));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R0_INV_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3398));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R1_INV_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R2_INV_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R2_INV_1 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3434));
  sky130_fd_sc_hd__clkbuf_4 T14Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3470));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R0_INV_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3506));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R1_INV_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R2_INV_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R2_INV_1 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3542));
  sky130_fd_sc_hd__clkbuf_4 T14Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3578));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R0_INV_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3614));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R1_INV_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R2_INV_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R2_INV_1 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3650));
  sky130_fd_sc_hd__clkbuf_4 T14Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3686));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R0_INV_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3722));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R1_INV_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R2_INV_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R2_INV_1 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3758));
  sky130_fd_sc_hd__clkbuf_4 T14Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3794));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R0_INV_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3830));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R1_INV_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R2_INV_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R2_INV_1 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3866));
  sky130_fd_sc_hd__clkbuf_4 T14Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3902));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R0_INV_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3938));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R1_INV_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R2_INV_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R2_INV_1 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3974));
  sky130_fd_sc_hd__clkbuf_4 T14Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4010));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R0_INV_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4046));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R1_INV_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R2_INV_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R2_INV_1 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4082));
  sky130_fd_sc_hd__clkbuf_4 T14Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4118));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R0_INV_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4154));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R1_INV_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R2_INV_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R2_INV_1 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4190));
  sky130_fd_sc_hd__clkbuf_4 T14Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4226));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R0_INV_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4262));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R1_INV_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R2_INV_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R2_INV_1 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4298));
  sky130_fd_sc_hd__clkbuf_4 T14Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B340));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R0_INV_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B375));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R1_INV_0 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R2_INV_0 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R2_INV_1 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B411));
  sky130_fd_sc_hd__clkbuf_4 T14Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4334));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R0_INV_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4370));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R1_INV_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R2_INV_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R2_INV_1 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4406));
  sky130_fd_sc_hd__clkbuf_4 T14Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4442));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R0_INV_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4478));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R1_INV_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R2_INV_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R2_INV_1 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4514));
  sky130_fd_sc_hd__clkbuf_4 T14Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4550));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R0_INV_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4586));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R1_INV_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R2_INV_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R2_INV_1 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4622));
  sky130_fd_sc_hd__clkbuf_4 T14Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4658));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R0_INV_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4694));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R1_INV_0 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R2_INV_0 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R2_INV_1 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4730));
  sky130_fd_sc_hd__clkbuf_4 T14Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4766));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R0_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4802));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R1_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R2_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R2_INV_1 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4838));
  sky130_fd_sc_hd__clkbuf_4 T14Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4874));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R0_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4910));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R1_INV_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R2_INV_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R2_INV_1 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4946));
  sky130_fd_sc_hd__clkbuf_4 T14Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4982));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R0_INV_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5018));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R1_INV_0 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R2_INV_0 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R2_INV_1 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5054));
  sky130_fd_sc_hd__clkbuf_4 T14Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5090));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R0_INV_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5126));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R1_INV_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R2_INV_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R2_INV_1 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5162));
  sky130_fd_sc_hd__clkbuf_4 T14Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5198));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R0_INV_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5234));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R1_INV_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R2_INV_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R2_INV_1 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5270));
  sky130_fd_sc_hd__clkbuf_4 T14Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5306));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R0_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5342));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R1_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R2_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R2_INV_1 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5378));
  sky130_fd_sc_hd__clkbuf_4 T14Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B447));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R0_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B483));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R1_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R2_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R2_INV_1 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B519));
  sky130_fd_sc_hd__clkbuf_4 T14Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5414));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R0_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5450));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R1_INV_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R2_INV_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R2_INV_1 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5486));
  sky130_fd_sc_hd__clkbuf_4 T14Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5522));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R0_INV_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5558));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R1_INV_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R2_INV_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R2_INV_1 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5594));
  sky130_fd_sc_hd__clkbuf_4 T14Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5630));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R0_INV_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5666));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R1_INV_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R2_INV_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R2_INV_1 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5702));
  sky130_fd_sc_hd__clkbuf_4 T14Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5738));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R0_INV_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5774));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R1_INV_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R2_INV_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R2_INV_1 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5810));
  sky130_fd_sc_hd__clkbuf_4 T14Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5846));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R0_INV_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5882));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R1_INV_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R2_INV_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R2_INV_1 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5918));
  sky130_fd_sc_hd__clkbuf_4 T14Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5954));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R0_INV_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5990));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R1_INV_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R2_INV_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R2_INV_1 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6026));
  sky130_fd_sc_hd__clkbuf_4 T14Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6062));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R0_INV_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6098));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R1_INV_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R2_INV_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R2_INV_1 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6134));
  sky130_fd_sc_hd__clkbuf_4 T14Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6170));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R0_INV_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6206));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R1_INV_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R2_INV_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R2_INV_1 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6242));
  sky130_fd_sc_hd__clkbuf_4 T14Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6278));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R0_INV_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6314));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R1_INV_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R2_INV_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R2_INV_1 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6350));
  sky130_fd_sc_hd__clkbuf_4 T14Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6386));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R0_INV_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6422));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R1_INV_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R2_INV_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R2_INV_1 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6458));
  sky130_fd_sc_hd__clkbuf_4 T14Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B555));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R0_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B591));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R1_INV_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R2_INV_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R2_INV_1 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B627));
  sky130_fd_sc_hd__clkbuf_4 T14Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6494));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R0_INV_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6530));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R1_INV_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R2_INV_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R2_INV_1 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6566));
  sky130_fd_sc_hd__clkbuf_4 T14Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6602));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R0_INV_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6638));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R1_INV_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R2_INV_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R2_INV_1 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6674));
  sky130_fd_sc_hd__clkbuf_4 T14Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6710));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R0_INV_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6746));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R1_INV_0 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R2_INV_0 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R2_INV_1 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6782));
  sky130_fd_sc_hd__clkbuf_4 T14Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6818));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R0_INV_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6854));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R1_INV_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R2_INV_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R2_INV_1 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6890));
  sky130_fd_sc_hd__clkbuf_4 T14Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6926));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R0_INV_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6962));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R1_INV_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R2_INV_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R2_INV_1 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6998));
  sky130_fd_sc_hd__clkbuf_4 T14Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7034));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R0_INV_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7070));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R1_INV_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R2_INV_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R2_INV_1 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7106));
  sky130_fd_sc_hd__clkbuf_4 T14Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7142));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R0_INV_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7178));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R1_INV_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R2_INV_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R2_INV_1 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7214));
  sky130_fd_sc_hd__clkbuf_4 T14Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7250));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R0_INV_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7286));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R1_INV_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R2_INV_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R2_INV_1 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7322));
  sky130_fd_sc_hd__clkbuf_4 T14Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7358));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R0_INV_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7394));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R1_INV_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R2_INV_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R2_INV_1 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7430));
  sky130_fd_sc_hd__clkbuf_4 T14Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7466));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R0_INV_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7502));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R1_INV_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R2_INV_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R2_INV_1 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7538));
  sky130_fd_sc_hd__clkbuf_4 T14Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B663));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R0_INV_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B699));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R1_INV_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R2_INV_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R2_INV_1 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B735));
  sky130_fd_sc_hd__clkbuf_4 T14Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7574));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R0_INV_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7610));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R1_INV_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R2_INV_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R2_INV_1 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7646));
  sky130_fd_sc_hd__clkbuf_4 T14Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7682));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R0_INV_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7718));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R1_INV_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R2_INV_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R2_INV_1 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7754));
  sky130_fd_sc_hd__clkbuf_4 T14Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7790));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R0_INV_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7826));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R1_INV_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R2_INV_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R2_INV_1 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7862));
  sky130_fd_sc_hd__clkbuf_4 T14Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7898));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R0_INV_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7934));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R1_INV_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R2_INV_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R2_INV_1 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7970));
  sky130_fd_sc_hd__clkbuf_4 T14Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8006));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R0_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8042));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R1_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R2_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R2_INV_1 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8078));
  sky130_fd_sc_hd__clkbuf_4 T14Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8114));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R0_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8150));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R1_INV_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R2_INV_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R2_INV_1 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8186));
  sky130_fd_sc_hd__clkbuf_4 T14Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8222));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R0_INV_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8258));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R1_INV_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R2_INV_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R2_INV_1 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8294));
  sky130_fd_sc_hd__clkbuf_4 T14Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8330));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R0_INV_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8366));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R1_INV_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R2_INV_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R2_INV_1 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8402));
  sky130_fd_sc_hd__clkbuf_4 T14Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8438));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R0_INV_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8474));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R1_INV_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R2_INV_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R2_INV_1 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8510));
  sky130_fd_sc_hd__clkbuf_4 T14Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8546));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R0_INV_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8582));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R1_INV_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R2_INV_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R2_INV_1 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8618));
  sky130_fd_sc_hd__clkbuf_4 T14Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B771));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R0_INV_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B807));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R1_INV_0 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R2_INV_0 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R2_INV_1 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B843));
  sky130_fd_sc_hd__clkbuf_4 T14Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8654));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R0_INV_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8690));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R1_INV_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R2_INV_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R2_INV_1 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8726));
  sky130_fd_sc_hd__clkbuf_4 T14Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8762));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R0_INV_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8798));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R1_INV_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R2_INV_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R2_INV_1 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8834));
  sky130_fd_sc_hd__clkbuf_4 T14Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8870));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R0_INV_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8906));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R1_INV_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R2_INV_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R2_INV_1 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8942));
  sky130_fd_sc_hd__clkbuf_4 T14Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8978));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R0_INV_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9014));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R1_INV_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R2_INV_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R2_INV_1 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9050));
  sky130_fd_sc_hd__clkbuf_4 T14Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9086));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R0_INV_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9122));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R1_INV_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R2_INV_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R2_INV_1 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9158));
  sky130_fd_sc_hd__clkbuf_4 T14Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9194));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R0_INV_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9230));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R1_INV_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R2_INV_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R2_INV_1 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9266));
  sky130_fd_sc_hd__clkbuf_4 T14Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9302));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R0_INV_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9338));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R1_INV_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R2_INV_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R2_INV_1 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9374));
  sky130_fd_sc_hd__clkbuf_4 T14Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9410));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R0_INV_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9446));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R1_INV_0 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R2_INV_0 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R2_INV_1 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9482));
  sky130_fd_sc_hd__clkbuf_4 T14Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9518));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R0_INV_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9554));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R1_INV_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R2_INV_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R2_INV_1 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9590));
  sky130_fd_sc_hd__clkbuf_4 T14Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9626));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R0_INV_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9662));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R1_INV_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R2_INV_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R2_INV_1 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9698));
  sky130_fd_sc_hd__clkbuf_4 T14Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B879));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R0_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B915));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R1_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R2_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R2_INV_1 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B951));
  sky130_fd_sc_hd__clkbuf_4 T14Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B987));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R0_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1023));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R1_INV_0 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R2_INV_0 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R2_INV_1 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1059));
  sky130_fd_sc_hd__clkbuf_4 T15Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B25));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R0_INV_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B60));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R1_INV_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R2_INV_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R2_INV_1 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B95));
  sky130_fd_sc_hd__clkbuf_4 T15Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1096));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R0_INV_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1132));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R1_INV_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R2_INV_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R2_INV_1 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y10__R3_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B73));
  sky130_fd_sc_hd__clkbuf_4 T15Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1204));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R0_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1240));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R1_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R2_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R2_INV_1 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1276));
  sky130_fd_sc_hd__clkbuf_4 T15Y12__R0_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B82));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R0_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1348));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R1_INV_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R2_INV_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R2_INV_1 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1384));
  sky130_fd_sc_hd__clkbuf_4 T15Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1420));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R0_INV_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y13__R1_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B91));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R1_INV_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R2_INV_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R2_INV_1 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1492));
  sky130_fd_sc_hd__clkbuf_4 T15Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1528));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R0_INV_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1563));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R1_INV_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R2_INV_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R2_INV_1 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1599));
  sky130_fd_sc_hd__clkbuf_4 T15Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1635));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R0_INV_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1671));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R1_INV_0 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R2_INV_0 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R2_INV_1 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1707));
  sky130_fd_sc_hd__clkbuf_4 T15Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1743));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R0_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1779));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R1_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R2_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R2_INV_1 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1815));
  sky130_fd_sc_hd__clkbuf_4 T15Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1851));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R0_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1887));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R1_INV_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R2_INV_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R2_INV_1 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1923));
  sky130_fd_sc_hd__clkbuf_4 T15Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1959));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R0_INV_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1995));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R1_INV_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R2_INV_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R2_INV_1 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2031));
  sky130_fd_sc_hd__clkbuf_4 T15Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2067));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R0_INV_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2103));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R1_INV_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R2_INV_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R2_INV_1 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2139));
  sky130_fd_sc_hd__clkbuf_4 T15Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B130));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R0_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B165));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R1_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R2_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R2_INV_1 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B200));
  sky130_fd_sc_hd__clkbuf_4 T15Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2175));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R0_INV_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2211));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R1_INV_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R2_INV_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R2_INV_1 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2247));
  sky130_fd_sc_hd__clkbuf_4 T15Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2283));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R0_INV_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2319));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R1_INV_0 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R2_INV_0 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R2_INV_1 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2355));
  sky130_fd_sc_hd__clkbuf_4 T15Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2391));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R0_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2427));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R1_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R2_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R2_INV_1 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2463));
  sky130_fd_sc_hd__clkbuf_4 T15Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2499));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R0_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2535));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R1_INV_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R2_INV_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R2_INV_1 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2571));
  sky130_fd_sc_hd__clkbuf_4 T15Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2607));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R0_INV_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2643));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R1_INV_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R2_INV_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R2_INV_1 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2679));
  sky130_fd_sc_hd__clkbuf_4 T15Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2715));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R0_INV_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2751));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R1_INV_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R2_INV_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R2_INV_1 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2787));
  sky130_fd_sc_hd__clkbuf_4 T15Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2823));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R0_INV_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2859));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R1_INV_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R2_INV_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R2_INV_1 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2895));
  sky130_fd_sc_hd__clkbuf_4 T15Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2931));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R0_INV_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2967));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R1_INV_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R2_INV_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R2_INV_1 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3003));
  sky130_fd_sc_hd__clkbuf_4 T15Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3039));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R0_INV_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3075));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R1_INV_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R2_INV_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R2_INV_1 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3111));
  sky130_fd_sc_hd__clkbuf_4 T15Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3147));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R0_INV_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3183));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R1_INV_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R2_INV_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R2_INV_1 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3219));
  sky130_fd_sc_hd__clkbuf_4 T15Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B235));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R0_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B270));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R1_INV_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R2_INV_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R2_INV_1 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B306));
  sky130_fd_sc_hd__clkbuf_4 T15Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3255));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R0_INV_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3291));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R1_INV_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R2_INV_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R2_INV_1 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3327));
  sky130_fd_sc_hd__clkbuf_4 T15Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3363));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R0_INV_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3399));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R1_INV_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R2_INV_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R2_INV_1 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3435));
  sky130_fd_sc_hd__clkbuf_4 T15Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3471));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R0_INV_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3507));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R1_INV_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R2_INV_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R2_INV_1 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3543));
  sky130_fd_sc_hd__clkbuf_4 T15Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3579));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R0_INV_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3615));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R1_INV_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R2_INV_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R2_INV_1 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3651));
  sky130_fd_sc_hd__clkbuf_4 T15Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3687));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R0_INV_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3723));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R1_INV_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R2_INV_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R2_INV_1 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3759));
  sky130_fd_sc_hd__clkbuf_4 T15Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3795));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R0_INV_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3831));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R1_INV_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R2_INV_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R2_INV_1 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3867));
  sky130_fd_sc_hd__clkbuf_4 T15Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3903));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R0_INV_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3939));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R1_INV_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R2_INV_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R2_INV_1 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3975));
  sky130_fd_sc_hd__clkbuf_4 T15Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4011));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R0_INV_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4047));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R1_INV_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R2_INV_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R2_INV_1 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4083));
  sky130_fd_sc_hd__clkbuf_4 T15Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4119));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R0_INV_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4155));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R1_INV_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R2_INV_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R2_INV_1 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4191));
  sky130_fd_sc_hd__clkbuf_4 T15Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4227));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R0_INV_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4263));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R1_INV_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R2_INV_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R2_INV_1 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4299));
  sky130_fd_sc_hd__clkbuf_4 T15Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B341));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R0_INV_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B376));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R1_INV_0 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R2_INV_0 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R2_INV_1 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B412));
  sky130_fd_sc_hd__clkbuf_4 T15Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4335));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R0_INV_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4371));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R1_INV_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R2_INV_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R2_INV_1 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4407));
  sky130_fd_sc_hd__clkbuf_4 T15Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4443));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R0_INV_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4479));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R1_INV_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R2_INV_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R2_INV_1 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4515));
  sky130_fd_sc_hd__clkbuf_4 T15Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4551));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R0_INV_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4587));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R1_INV_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R2_INV_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R2_INV_1 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4623));
  sky130_fd_sc_hd__clkbuf_4 T15Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4659));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R0_INV_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4695));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R1_INV_0 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R2_INV_0 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R2_INV_1 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4731));
  sky130_fd_sc_hd__clkbuf_4 T15Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4767));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R0_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4803));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R1_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R2_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R2_INV_1 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4839));
  sky130_fd_sc_hd__clkbuf_4 T15Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4875));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R0_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4911));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R1_INV_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R2_INV_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R2_INV_1 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4947));
  sky130_fd_sc_hd__clkbuf_4 T15Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4983));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R0_INV_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5019));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R1_INV_0 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R2_INV_0 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R2_INV_1 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5055));
  sky130_fd_sc_hd__clkbuf_4 T15Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5091));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R0_INV_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5127));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R1_INV_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R2_INV_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R2_INV_1 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5163));
  sky130_fd_sc_hd__clkbuf_4 T15Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5199));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R0_INV_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5235));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R1_INV_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R2_INV_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R2_INV_1 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5271));
  sky130_fd_sc_hd__clkbuf_4 T15Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5307));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R0_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5343));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R1_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R2_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R2_INV_1 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5379));
  sky130_fd_sc_hd__clkbuf_4 T15Y4__R0_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B28));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R0_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B484));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R1_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R2_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R2_INV_1 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B520));
  sky130_fd_sc_hd__clkbuf_4 T15Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5415));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R0_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5451));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R1_INV_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R2_INV_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R2_INV_1 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5487));
  sky130_fd_sc_hd__clkbuf_4 T15Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5523));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R0_INV_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5559));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R1_INV_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R2_INV_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R2_INV_1 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5595));
  sky130_fd_sc_hd__clkbuf_4 T15Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5631));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R0_INV_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5667));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R1_INV_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R2_INV_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R2_INV_1 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5703));
  sky130_fd_sc_hd__clkbuf_4 T15Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5739));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R0_INV_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5775));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R1_INV_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R2_INV_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R2_INV_1 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5811));
  sky130_fd_sc_hd__clkbuf_4 T15Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5847));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R0_INV_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5883));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R1_INV_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R2_INV_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R2_INV_1 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5919));
  sky130_fd_sc_hd__clkbuf_4 T15Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5955));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R0_INV_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5991));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R1_INV_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R2_INV_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R2_INV_1 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6027));
  sky130_fd_sc_hd__clkbuf_4 T15Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6063));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R0_INV_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6099));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R1_INV_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R2_INV_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R2_INV_1 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6135));
  sky130_fd_sc_hd__clkbuf_4 T15Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6171));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R0_INV_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6207));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R1_INV_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R2_INV_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R2_INV_1 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6243));
  sky130_fd_sc_hd__clkbuf_4 T15Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6279));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R0_INV_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6315));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R1_INV_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R2_INV_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R2_INV_1 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6351));
  sky130_fd_sc_hd__clkbuf_4 T15Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6387));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R0_INV_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6423));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R1_INV_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R2_INV_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R2_INV_1 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6459));
  sky130_fd_sc_hd__clkbuf_4 T15Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B556));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R0_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y5__R1_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B37));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R1_INV_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R2_INV_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R2_INV_1 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B628));
  sky130_fd_sc_hd__clkbuf_4 T15Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6495));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R0_INV_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6531));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R1_INV_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R2_INV_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R2_INV_1 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6567));
  sky130_fd_sc_hd__clkbuf_4 T15Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6603));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R0_INV_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6639));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R1_INV_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R2_INV_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R2_INV_1 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6675));
  sky130_fd_sc_hd__clkbuf_4 T15Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6711));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R0_INV_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6747));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R1_INV_0 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R2_INV_0 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R2_INV_1 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6783));
  sky130_fd_sc_hd__clkbuf_4 T15Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6819));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R0_INV_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6855));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R1_INV_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R2_INV_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R2_INV_1 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6891));
  sky130_fd_sc_hd__clkbuf_4 T15Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6927));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R0_INV_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6963));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R1_INV_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R2_INV_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R2_INV_1 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6999));
  sky130_fd_sc_hd__clkbuf_4 T15Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7035));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R0_INV_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7071));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R1_INV_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R2_INV_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R2_INV_1 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7107));
  sky130_fd_sc_hd__clkbuf_4 T15Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7143));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R0_INV_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7179));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R1_INV_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R2_INV_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R2_INV_1 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7215));
  sky130_fd_sc_hd__clkbuf_4 T15Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7251));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R0_INV_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7287));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R1_INV_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R2_INV_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R2_INV_1 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7323));
  sky130_fd_sc_hd__clkbuf_4 T15Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7359));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R0_INV_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7395));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R1_INV_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R2_INV_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R2_INV_1 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7431));
  sky130_fd_sc_hd__clkbuf_4 T15Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7467));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R0_INV_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7503));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R1_INV_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R2_INV_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R2_INV_1 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7539));
  sky130_fd_sc_hd__clkbuf_4 T15Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B664));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R0_INV_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B700));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R1_INV_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R2_INV_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R2_INV_1 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y6__R3_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B46));
  sky130_fd_sc_hd__clkbuf_4 T15Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7575));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R0_INV_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7611));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R1_INV_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R2_INV_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R2_INV_1 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7647));
  sky130_fd_sc_hd__clkbuf_4 T15Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7683));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R0_INV_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7719));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R1_INV_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R2_INV_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R2_INV_1 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7755));
  sky130_fd_sc_hd__clkbuf_4 T15Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7791));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R0_INV_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7827));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R1_INV_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R2_INV_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R2_INV_1 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7863));
  sky130_fd_sc_hd__clkbuf_4 T15Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7899));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R0_INV_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7935));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R1_INV_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R2_INV_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R2_INV_1 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7971));
  sky130_fd_sc_hd__clkbuf_4 T15Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8007));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R0_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8043));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R1_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R2_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R2_INV_1 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8079));
  sky130_fd_sc_hd__clkbuf_4 T15Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8115));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R0_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8151));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R1_INV_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R2_INV_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R2_INV_1 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8187));
  sky130_fd_sc_hd__clkbuf_4 T15Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8223));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R0_INV_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8259));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R1_INV_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R2_INV_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R2_INV_1 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8295));
  sky130_fd_sc_hd__clkbuf_4 T15Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8331));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R0_INV_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8367));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R1_INV_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R2_INV_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R2_INV_1 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8403));
  sky130_fd_sc_hd__clkbuf_4 T15Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8439));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R0_INV_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8475));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R1_INV_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R2_INV_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R2_INV_1 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8511));
  sky130_fd_sc_hd__clkbuf_4 T15Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8547));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R0_INV_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8583));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R1_INV_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R2_INV_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R2_INV_1 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8619));
  sky130_fd_sc_hd__clkbuf_4 T15Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B772));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R0_INV_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B808));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R1_INV_0 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R2_INV_0 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R2_INV_1 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B844));
  sky130_fd_sc_hd__clkbuf_4 T15Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8655));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R0_INV_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8691));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R1_INV_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R2_INV_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R2_INV_1 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8727));
  sky130_fd_sc_hd__clkbuf_4 T15Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8763));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R0_INV_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8799));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R1_INV_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R2_INV_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R2_INV_1 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8835));
  sky130_fd_sc_hd__clkbuf_4 T15Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8871));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R0_INV_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8907));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R1_INV_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R2_INV_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R2_INV_1 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8943));
  sky130_fd_sc_hd__clkbuf_4 T15Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8979));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R0_INV_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9015));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R1_INV_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R2_INV_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R2_INV_1 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9051));
  sky130_fd_sc_hd__clkbuf_4 T15Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9087));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R0_INV_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9123));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R1_INV_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R2_INV_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R2_INV_1 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9159));
  sky130_fd_sc_hd__clkbuf_4 T15Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9195));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R0_INV_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9231));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R1_INV_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R2_INV_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R2_INV_1 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9267));
  sky130_fd_sc_hd__clkbuf_4 T15Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9303));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R0_INV_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9339));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R1_INV_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R2_INV_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R2_INV_1 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9375));
  sky130_fd_sc_hd__clkbuf_4 T15Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9411));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R0_INV_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9447));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R1_INV_0 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R2_INV_0 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R2_INV_1 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9483));
  sky130_fd_sc_hd__clkbuf_4 T15Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9519));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R0_INV_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9555));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R1_INV_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R2_INV_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R2_INV_1 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9591));
  sky130_fd_sc_hd__clkbuf_4 T15Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9627));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R0_INV_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9663));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R1_INV_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R2_INV_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R2_INV_1 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9699));
  sky130_fd_sc_hd__clkbuf_4 T15Y8__R0_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B55));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R0_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B916));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R1_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R2_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R2_INV_1 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B952));
  sky130_fd_sc_hd__clkbuf_4 T15Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B988));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R0_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y9__R1_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B4));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R1_INV_0 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R2_INV_0 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R2_INV_1 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1060));
  sky130_fd_sc_hd__clkbuf_4 T16Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B26));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R0_INV_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B61));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R1_INV_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R2_INV_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R2_INV_1 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y0__R3_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B6));
  sky130_fd_sc_hd__clkbuf_4 T16Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1097));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R0_INV_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1133));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R1_INV_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R2_INV_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R2_INV_1 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1169));
  sky130_fd_sc_hd__clkbuf_4 T16Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1205));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R0_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1241));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R1_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R2_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R2_INV_1 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1277));
  sky130_fd_sc_hd__clkbuf_4 T16Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1313));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R0_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1349));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R1_INV_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R2_INV_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R2_INV_1 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1385));
  sky130_fd_sc_hd__clkbuf_4 T16Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1421));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R0_INV_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1457));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R1_INV_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R2_INV_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R2_INV_1 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1493));
  sky130_fd_sc_hd__clkbuf_4 T16Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1529));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R0_INV_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1564));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R1_INV_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R2_INV_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R2_INV_1 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y14__R3_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B100));
  sky130_fd_sc_hd__clkbuf_4 T16Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1636));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R0_INV_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1672));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R1_INV_0 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R2_INV_0 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R2_INV_1 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1708));
  sky130_fd_sc_hd__clkbuf_4 T16Y16__R0_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B109));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R0_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1780));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R1_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R2_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R2_INV_1 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1816));
  sky130_fd_sc_hd__clkbuf_4 T16Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1852));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R0_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y17__R1_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B118));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R1_INV_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R2_INV_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R2_INV_1 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1924));
  sky130_fd_sc_hd__clkbuf_4 T16Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1960));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R0_INV_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1996));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R1_INV_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R2_INV_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R2_INV_1 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y18__R3_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B127));
  sky130_fd_sc_hd__clkbuf_4 T16Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2068));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R0_INV_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2104));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R1_INV_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R2_INV_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R2_INV_1 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2140));
  sky130_fd_sc_hd__clkbuf_4 T16Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B131));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R0_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B166));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R1_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R2_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R2_INV_1 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B201));
  sky130_fd_sc_hd__clkbuf_4 T16Y20__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B136));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R0_INV_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2212));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R1_INV_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R2_INV_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R2_INV_1 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2248));
  sky130_fd_sc_hd__clkbuf_4 T16Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2284));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R0_INV_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y21__R1_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B145));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R1_INV_0 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R2_INV_0 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R2_INV_1 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2356));
  sky130_fd_sc_hd__clkbuf_4 T16Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2392));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R0_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2428));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R1_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R2_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R2_INV_1 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y22__R3_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B154));
  sky130_fd_sc_hd__clkbuf_4 T16Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2500));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R0_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2536));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R1_INV_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R2_INV_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R2_INV_1 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2572));
  sky130_fd_sc_hd__clkbuf_4 T16Y24__R0_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B163));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R0_INV_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2644));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R1_INV_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R2_INV_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R2_INV_1 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2680));
  sky130_fd_sc_hd__clkbuf_4 T16Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2716));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R0_INV_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y25__R1_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B172));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R1_INV_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R2_INV_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R2_INV_1 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2788));
  sky130_fd_sc_hd__clkbuf_4 T16Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2824));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R0_INV_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2860));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R1_INV_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R2_INV_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R2_INV_1 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y26__R3_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B181));
  sky130_fd_sc_hd__clkbuf_4 T16Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2932));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R0_INV_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2968));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R1_INV_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R2_INV_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R2_INV_1 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3004));
  sky130_fd_sc_hd__clkbuf_4 T16Y28__R0_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B190));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R0_INV_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3076));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R1_INV_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R2_INV_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R2_INV_1 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3112));
  sky130_fd_sc_hd__clkbuf_4 T16Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3148));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R0_INV_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y29__R1_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B199));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R1_INV_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R2_INV_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R2_INV_1 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3220));
  sky130_fd_sc_hd__clkbuf_4 T16Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B236));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R0_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B271));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R1_INV_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R2_INV_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R2_INV_1 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B307));
  sky130_fd_sc_hd__clkbuf_4 T16Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3256));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R0_INV_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3292));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R1_INV_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R2_INV_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R2_INV_1 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y30__R3_BUF_0 (.A(clk_L4_B0), .X(clk_L3_B1));
  sky130_fd_sc_hd__clkbuf_4 T16Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3364));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R0_INV_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3400));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R1_INV_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R2_INV_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R2_INV_1 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3436));
  sky130_fd_sc_hd__clkbuf_4 T16Y32__R0_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B217));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R0_INV_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3508));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R1_INV_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R2_INV_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R2_INV_1 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3544));
  sky130_fd_sc_hd__clkbuf_4 T16Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3580));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R0_INV_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y33__R1_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B226));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R1_INV_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R2_INV_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R2_INV_1 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3652));
  sky130_fd_sc_hd__clkbuf_4 T16Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3688));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R0_INV_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3724));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R1_INV_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R2_INV_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R2_INV_1 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y34__R3_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B235));
  sky130_fd_sc_hd__clkbuf_4 T16Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3796));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R0_INV_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3832));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R1_INV_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R2_INV_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R2_INV_1 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3868));
  sky130_fd_sc_hd__clkbuf_4 T16Y36__R0_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B244));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R0_INV_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3940));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R1_INV_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R2_INV_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R2_INV_1 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3976));
  sky130_fd_sc_hd__clkbuf_4 T16Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4012));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R0_INV_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y37__R1_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B253));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R1_INV_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R2_INV_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R2_INV_1 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4084));
  sky130_fd_sc_hd__clkbuf_4 T16Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4120));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R0_INV_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4156));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R1_INV_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R2_INV_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R2_INV_1 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y38__R3_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B262));
  sky130_fd_sc_hd__clkbuf_4 T16Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4228));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R0_INV_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4264));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R1_INV_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R2_INV_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R2_INV_1 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4300));
  sky130_fd_sc_hd__clkbuf_4 T16Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B342));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R0_INV_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B377));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R1_INV_0 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R2_INV_0 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R2_INV_1 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B413));
  sky130_fd_sc_hd__clkbuf_4 T16Y40__R0_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B271));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R0_INV_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4372));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R1_INV_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R2_INV_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R2_INV_1 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4408));
  sky130_fd_sc_hd__clkbuf_4 T16Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4444));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R0_INV_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y41__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B280));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R1_INV_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R2_INV_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R2_INV_1 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4516));
  sky130_fd_sc_hd__clkbuf_4 T16Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4552));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R0_INV_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4588));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R1_INV_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R2_INV_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R2_INV_1 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y42__R3_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B289));
  sky130_fd_sc_hd__clkbuf_4 T16Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4660));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R0_INV_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4696));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R1_INV_0 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R2_INV_0 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R2_INV_1 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4732));
  sky130_fd_sc_hd__clkbuf_4 T16Y44__R0_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B298));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R0_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4804));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R1_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R2_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R2_INV_1 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4840));
  sky130_fd_sc_hd__clkbuf_4 T16Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4876));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R0_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y45__R1_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B307));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R1_INV_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R2_INV_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R2_INV_1 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4948));
  sky130_fd_sc_hd__clkbuf_4 T16Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4984));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R0_INV_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5020));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R1_INV_0 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R2_INV_0 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R2_INV_1 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y46__R3_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B316));
  sky130_fd_sc_hd__clkbuf_4 T16Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5092));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R0_INV_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5128));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R1_INV_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R2_INV_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R2_INV_1 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5164));
  sky130_fd_sc_hd__clkbuf_4 T16Y48__R0_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B325));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R0_INV_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5236));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R1_INV_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R2_INV_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R2_INV_1 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5272));
  sky130_fd_sc_hd__clkbuf_4 T16Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5308));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R0_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y49__R1_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B334));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R1_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R2_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R2_INV_1 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5380));
  sky130_fd_sc_hd__clkbuf_4 T16Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B449));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R0_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B485));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R1_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R2_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R2_INV_1 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B521));
  sky130_fd_sc_hd__clkbuf_4 T16Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5416));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R0_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5452));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R1_INV_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R2_INV_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R2_INV_1 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y50__R3_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B343));
  sky130_fd_sc_hd__clkbuf_4 T16Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5524));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R0_INV_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5560));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R1_INV_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R2_INV_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R2_INV_1 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5596));
  sky130_fd_sc_hd__clkbuf_4 T16Y52__R0_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B22));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R0_INV_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5668));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R1_INV_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R2_INV_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R2_INV_1 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5704));
  sky130_fd_sc_hd__clkbuf_4 T16Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5740));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R0_INV_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y53__R1_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B361));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R1_INV_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R2_INV_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R2_INV_1 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5812));
  sky130_fd_sc_hd__clkbuf_4 T16Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5848));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R0_INV_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5884));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R1_INV_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R2_INV_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R2_INV_1 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y54__R3_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B370));
  sky130_fd_sc_hd__clkbuf_4 T16Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5956));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R0_INV_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5992));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R1_INV_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R2_INV_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R2_INV_1 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6028));
  sky130_fd_sc_hd__clkbuf_4 T16Y56__R0_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B379));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R0_INV_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6100));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R1_INV_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R2_INV_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R2_INV_1 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6136));
  sky130_fd_sc_hd__clkbuf_4 T16Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6172));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R0_INV_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y57__R1_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B388));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R1_INV_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R2_INV_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R2_INV_1 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6244));
  sky130_fd_sc_hd__clkbuf_4 T16Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6280));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R0_INV_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6316));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R1_INV_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R2_INV_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R2_INV_1 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y58__R3_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B397));
  sky130_fd_sc_hd__clkbuf_4 T16Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6388));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R0_INV_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6424));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R1_INV_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R2_INV_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R2_INV_1 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6460));
  sky130_fd_sc_hd__clkbuf_4 T16Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B557));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R0_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B593));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R1_INV_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R2_INV_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R2_INV_1 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B629));
  sky130_fd_sc_hd__clkbuf_4 T16Y60__R0_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B406));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R0_INV_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6532));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R1_INV_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R2_INV_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R2_INV_1 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6568));
  sky130_fd_sc_hd__clkbuf_4 T16Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6604));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R0_INV_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y61__R1_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B415));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R1_INV_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R2_INV_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R2_INV_1 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6676));
  sky130_fd_sc_hd__clkbuf_4 T16Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6712));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R0_INV_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6748));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R1_INV_0 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R2_INV_0 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R2_INV_1 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y62__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B424));
  sky130_fd_sc_hd__clkbuf_4 T16Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6820));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R0_INV_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6856));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R1_INV_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R2_INV_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R2_INV_1 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6892));
  sky130_fd_sc_hd__clkbuf_4 T16Y64__R0_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B433));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R0_INV_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6964));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R1_INV_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R2_INV_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R2_INV_1 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7000));
  sky130_fd_sc_hd__clkbuf_4 T16Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7036));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R0_INV_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y65__R1_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B442));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R1_INV_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R2_INV_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R2_INV_1 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7108));
  sky130_fd_sc_hd__clkbuf_4 T16Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7144));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R0_INV_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7180));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R1_INV_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R2_INV_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R2_INV_1 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y66__R3_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B451));
  sky130_fd_sc_hd__clkbuf_4 T16Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7252));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R0_INV_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7288));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R1_INV_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R2_INV_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R2_INV_1 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7324));
  sky130_fd_sc_hd__clkbuf_4 T16Y68__R0_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B460));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R0_INV_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7396));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R1_INV_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R2_INV_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R2_INV_1 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7432));
  sky130_fd_sc_hd__clkbuf_4 T16Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7468));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R0_INV_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y69__R1_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B469));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R1_INV_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R2_INV_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R2_INV_1 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7540));
  sky130_fd_sc_hd__clkbuf_4 T16Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B665));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R0_INV_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B701));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R1_INV_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R2_INV_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R2_INV_1 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B737));
  sky130_fd_sc_hd__clkbuf_4 T16Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7576));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R0_INV_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7612));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R1_INV_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R2_INV_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R2_INV_1 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y70__R3_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B478));
  sky130_fd_sc_hd__clkbuf_4 T16Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7684));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R0_INV_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7720));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R1_INV_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R2_INV_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R2_INV_1 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7756));
  sky130_fd_sc_hd__clkbuf_4 T16Y72__R0_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B487));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R0_INV_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7828));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R1_INV_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R2_INV_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R2_INV_1 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7864));
  sky130_fd_sc_hd__clkbuf_4 T16Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7900));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R0_INV_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y73__R1_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B31));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R1_INV_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R2_INV_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R2_INV_1 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7972));
  sky130_fd_sc_hd__clkbuf_4 T16Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8008));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R0_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8044));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R1_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R2_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R2_INV_1 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y74__R3_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B505));
  sky130_fd_sc_hd__clkbuf_4 T16Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8116));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R0_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8152));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R1_INV_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R2_INV_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R2_INV_1 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8188));
  sky130_fd_sc_hd__clkbuf_4 T16Y76__R0_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B514));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R0_INV_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8260));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R1_INV_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R2_INV_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R2_INV_1 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8296));
  sky130_fd_sc_hd__clkbuf_4 T16Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8332));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R0_INV_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y77__R1_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B523));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R1_INV_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R2_INV_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R2_INV_1 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8404));
  sky130_fd_sc_hd__clkbuf_4 T16Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8440));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R0_INV_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8476));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R1_INV_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R2_INV_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R2_INV_1 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y78__R3_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B532));
  sky130_fd_sc_hd__clkbuf_4 T16Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8548));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R0_INV_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8584));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R1_INV_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R2_INV_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R2_INV_1 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8620));
  sky130_fd_sc_hd__clkbuf_4 T16Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B773));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R0_INV_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B809));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R1_INV_0 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R2_INV_0 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R2_INV_1 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B845));
  sky130_fd_sc_hd__clkbuf_4 T16Y80__R0_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B541));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R0_INV_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8692));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R1_INV_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R2_INV_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R2_INV_1 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8728));
  sky130_fd_sc_hd__clkbuf_4 T16Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8764));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R0_INV_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y81__R1_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B550));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R1_INV_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R2_INV_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R2_INV_1 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8836));
  sky130_fd_sc_hd__clkbuf_4 T16Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8872));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R0_INV_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8908));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R1_INV_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R2_INV_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R2_INV_1 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y82__R3_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B559));
  sky130_fd_sc_hd__clkbuf_4 T16Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8980));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R0_INV_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9016));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R1_INV_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R2_INV_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R2_INV_1 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9052));
  sky130_fd_sc_hd__clkbuf_4 T16Y84__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B568));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R0_INV_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9124));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R1_INV_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R2_INV_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R2_INV_1 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9160));
  sky130_fd_sc_hd__clkbuf_4 T16Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9196));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R0_INV_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y85__R1_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B577));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R1_INV_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R2_INV_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R2_INV_1 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9268));
  sky130_fd_sc_hd__clkbuf_4 T16Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9304));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R0_INV_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9340));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R1_INV_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R2_INV_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R2_INV_1 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y86__R3_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B586));
  sky130_fd_sc_hd__clkbuf_4 T16Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9412));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R0_INV_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9448));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R1_INV_0 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R2_INV_0 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R2_INV_1 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9484));
  sky130_fd_sc_hd__clkbuf_4 T16Y88__R0_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B595));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R0_INV_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9556));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R1_INV_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R2_INV_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R2_INV_1 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9592));
  sky130_fd_sc_hd__clkbuf_4 T16Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9628));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R0_INV_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y89__R1_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B604));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R1_INV_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R2_INV_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R2_INV_1 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9700));
  sky130_fd_sc_hd__clkbuf_4 T16Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B881));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R0_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B917));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R1_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R2_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R2_INV_1 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B953));
  sky130_fd_sc_hd__clkbuf_4 T16Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B989));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R0_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1025));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R1_INV_0 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R2_INV_0 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R2_INV_1 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1061));
  sky130_fd_sc_hd__clkbuf_4 T17Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B27));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R0_INV_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B62));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R1_INV_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R2_INV_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R2_INV_1 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B97));
  sky130_fd_sc_hd__clkbuf_4 T17Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1098));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R0_INV_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1134));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R1_INV_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R2_INV_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R2_INV_1 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1170));
  sky130_fd_sc_hd__clkbuf_4 T17Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1206));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R0_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1242));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R1_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R2_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R2_INV_1 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1278));
  sky130_fd_sc_hd__clkbuf_4 T17Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1314));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R0_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1350));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R1_INV_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R2_INV_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R2_INV_1 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1386));
  sky130_fd_sc_hd__clkbuf_4 T17Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1422));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R0_INV_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1458));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R1_INV_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R2_INV_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R2_INV_1 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1494));
  sky130_fd_sc_hd__clkbuf_4 T17Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1530));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R0_INV_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1565));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R1_INV_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R2_INV_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R2_INV_1 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1601));
  sky130_fd_sc_hd__clkbuf_4 T17Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1637));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R0_INV_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1673));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R1_INV_0 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R2_INV_0 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R2_INV_1 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1709));
  sky130_fd_sc_hd__clkbuf_4 T17Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1745));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R0_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1781));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R1_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R2_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R2_INV_1 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1817));
  sky130_fd_sc_hd__clkbuf_4 T17Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1853));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R0_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1889));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R1_INV_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R2_INV_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R2_INV_1 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1925));
  sky130_fd_sc_hd__clkbuf_4 T17Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1961));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R0_INV_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1997));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R1_INV_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R2_INV_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R2_INV_1 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2033));
  sky130_fd_sc_hd__clkbuf_4 T17Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2069));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R0_INV_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2105));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R1_INV_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R2_INV_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R2_INV_1 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2141));
  sky130_fd_sc_hd__clkbuf_4 T17Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B132));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R0_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B167));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R1_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R2_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R2_INV_1 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B202));
  sky130_fd_sc_hd__clkbuf_4 T17Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2177));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R0_INV_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2213));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R1_INV_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R2_INV_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R2_INV_1 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2249));
  sky130_fd_sc_hd__clkbuf_4 T17Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2285));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R0_INV_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2321));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R1_INV_0 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R2_INV_0 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R2_INV_1 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2357));
  sky130_fd_sc_hd__clkbuf_4 T17Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2393));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R0_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2429));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R1_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R2_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R2_INV_1 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2465));
  sky130_fd_sc_hd__clkbuf_4 T17Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2501));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R0_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2537));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R1_INV_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R2_INV_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R2_INV_1 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2573));
  sky130_fd_sc_hd__clkbuf_4 T17Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2609));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R0_INV_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2645));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R1_INV_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R2_INV_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R2_INV_1 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2681));
  sky130_fd_sc_hd__clkbuf_4 T17Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2717));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R0_INV_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2753));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R1_INV_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R2_INV_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R2_INV_1 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2789));
  sky130_fd_sc_hd__clkbuf_4 T17Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2825));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R0_INV_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2861));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R1_INV_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R2_INV_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R2_INV_1 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2897));
  sky130_fd_sc_hd__clkbuf_4 T17Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2933));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R0_INV_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2969));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R1_INV_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R2_INV_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R2_INV_1 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3005));
  sky130_fd_sc_hd__clkbuf_4 T17Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3041));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R0_INV_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3077));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R1_INV_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R2_INV_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R2_INV_1 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3113));
  sky130_fd_sc_hd__clkbuf_4 T17Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3149));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R0_INV_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3185));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R1_INV_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R2_INV_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R2_INV_1 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3221));
  sky130_fd_sc_hd__clkbuf_4 T17Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B237));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R0_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y2__R1_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B17));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R1_INV_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R2_INV_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R2_INV_1 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B308));
  sky130_fd_sc_hd__clkbuf_4 T17Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3257));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R0_INV_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3293));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R1_INV_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R2_INV_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R2_INV_1 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3329));
  sky130_fd_sc_hd__clkbuf_4 T17Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3365));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R0_INV_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3401));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R1_INV_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R2_INV_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R2_INV_1 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3437));
  sky130_fd_sc_hd__clkbuf_4 T17Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3473));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R0_INV_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3509));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R1_INV_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R2_INV_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R2_INV_1 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3545));
  sky130_fd_sc_hd__clkbuf_4 T17Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3581));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R0_INV_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3617));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R1_INV_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R2_INV_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R2_INV_1 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3653));
  sky130_fd_sc_hd__clkbuf_4 T17Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3689));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R0_INV_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3725));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R1_INV_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R2_INV_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R2_INV_1 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3761));
  sky130_fd_sc_hd__clkbuf_4 T17Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3797));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R0_INV_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3833));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R1_INV_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R2_INV_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R2_INV_1 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3869));
  sky130_fd_sc_hd__clkbuf_4 T17Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3905));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R0_INV_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3941));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R1_INV_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R2_INV_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R2_INV_1 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3977));
  sky130_fd_sc_hd__clkbuf_4 T17Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4013));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R0_INV_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4049));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R1_INV_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R2_INV_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R2_INV_1 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4085));
  sky130_fd_sc_hd__clkbuf_4 T17Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4121));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R0_INV_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4157));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R1_INV_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R2_INV_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R2_INV_1 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4193));
  sky130_fd_sc_hd__clkbuf_4 T17Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4229));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R0_INV_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4265));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R1_INV_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R2_INV_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R2_INV_1 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4301));
  sky130_fd_sc_hd__clkbuf_4 T17Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B343));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R0_INV_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B378));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R1_INV_0 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R2_INV_0 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R2_INV_1 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B414));
  sky130_fd_sc_hd__clkbuf_4 T17Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4337));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R0_INV_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4373));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R1_INV_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R2_INV_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R2_INV_1 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4409));
  sky130_fd_sc_hd__clkbuf_4 T17Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4445));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R0_INV_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4481));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R1_INV_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R2_INV_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R2_INV_1 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4517));
  sky130_fd_sc_hd__clkbuf_4 T17Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4553));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R0_INV_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4589));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R1_INV_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R2_INV_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R2_INV_1 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4625));
  sky130_fd_sc_hd__clkbuf_4 T17Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4661));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R0_INV_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4697));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R1_INV_0 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R2_INV_0 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R2_INV_1 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4733));
  sky130_fd_sc_hd__clkbuf_4 T17Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4769));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R0_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4805));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R1_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R2_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R2_INV_1 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4841));
  sky130_fd_sc_hd__clkbuf_4 T17Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4877));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R0_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4913));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R1_INV_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R2_INV_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R2_INV_1 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4949));
  sky130_fd_sc_hd__clkbuf_4 T17Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4985));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R0_INV_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5021));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R1_INV_0 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R2_INV_0 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R2_INV_1 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5057));
  sky130_fd_sc_hd__clkbuf_4 T17Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5093));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R0_INV_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5129));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R1_INV_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R2_INV_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R2_INV_1 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5165));
  sky130_fd_sc_hd__clkbuf_4 T17Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5201));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R0_INV_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5237));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R1_INV_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R2_INV_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R2_INV_1 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5273));
  sky130_fd_sc_hd__clkbuf_4 T17Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5309));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R0_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5345));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R1_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R2_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R2_INV_1 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5381));
  sky130_fd_sc_hd__clkbuf_4 T17Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B450));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R0_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B486));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R1_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R2_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R2_INV_1 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B522));
  sky130_fd_sc_hd__clkbuf_4 T17Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5417));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R0_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5453));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R1_INV_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R2_INV_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R2_INV_1 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5489));
  sky130_fd_sc_hd__clkbuf_4 T17Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5525));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R0_INV_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5561));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R1_INV_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R2_INV_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R2_INV_1 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5597));
  sky130_fd_sc_hd__clkbuf_4 T17Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5633));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R0_INV_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5669));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R1_INV_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R2_INV_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R2_INV_1 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5705));
  sky130_fd_sc_hd__clkbuf_4 T17Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5741));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R0_INV_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5777));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R1_INV_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R2_INV_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R2_INV_1 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5813));
  sky130_fd_sc_hd__clkbuf_4 T17Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5849));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R0_INV_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5885));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R1_INV_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R2_INV_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R2_INV_1 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5921));
  sky130_fd_sc_hd__clkbuf_4 T17Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5957));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R0_INV_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5993));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R1_INV_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R2_INV_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R2_INV_1 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6029));
  sky130_fd_sc_hd__clkbuf_4 T17Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6065));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R0_INV_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6101));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R1_INV_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R2_INV_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R2_INV_1 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6137));
  sky130_fd_sc_hd__clkbuf_4 T17Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6173));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R0_INV_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6209));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R1_INV_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R2_INV_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R2_INV_1 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6245));
  sky130_fd_sc_hd__clkbuf_4 T17Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6281));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R0_INV_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6317));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R1_INV_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R2_INV_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R2_INV_1 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6353));
  sky130_fd_sc_hd__clkbuf_4 T17Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6389));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R0_INV_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6425));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R1_INV_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R2_INV_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R2_INV_1 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6461));
  sky130_fd_sc_hd__clkbuf_4 T17Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B558));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R0_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B594));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R1_INV_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R2_INV_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R2_INV_1 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B630));
  sky130_fd_sc_hd__clkbuf_4 T17Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6497));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R0_INV_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6533));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R1_INV_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R2_INV_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R2_INV_1 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6569));
  sky130_fd_sc_hd__clkbuf_4 T17Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6605));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R0_INV_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6641));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R1_INV_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R2_INV_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R2_INV_1 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6677));
  sky130_fd_sc_hd__clkbuf_4 T17Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6713));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R0_INV_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6749));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R1_INV_0 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R2_INV_0 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R2_INV_1 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6785));
  sky130_fd_sc_hd__clkbuf_4 T17Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6821));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R0_INV_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6857));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R1_INV_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R2_INV_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R2_INV_1 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6893));
  sky130_fd_sc_hd__clkbuf_4 T17Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6929));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R0_INV_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6965));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R1_INV_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R2_INV_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R2_INV_1 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7001));
  sky130_fd_sc_hd__clkbuf_4 T17Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7037));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R0_INV_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7073));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R1_INV_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R2_INV_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R2_INV_1 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7109));
  sky130_fd_sc_hd__clkbuf_4 T17Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7145));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R0_INV_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7181));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R1_INV_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R2_INV_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R2_INV_1 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7217));
  sky130_fd_sc_hd__clkbuf_4 T17Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7253));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R0_INV_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7289));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R1_INV_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R2_INV_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R2_INV_1 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7325));
  sky130_fd_sc_hd__clkbuf_4 T17Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7361));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R0_INV_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7397));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R1_INV_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R2_INV_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R2_INV_1 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7433));
  sky130_fd_sc_hd__clkbuf_4 T17Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7469));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R0_INV_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7505));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R1_INV_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R2_INV_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R2_INV_1 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7541));
  sky130_fd_sc_hd__clkbuf_4 T17Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B666));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R0_INV_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B702));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R1_INV_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R2_INV_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R2_INV_1 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B738));
  sky130_fd_sc_hd__clkbuf_4 T17Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7577));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R0_INV_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7613));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R1_INV_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R2_INV_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R2_INV_1 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7649));
  sky130_fd_sc_hd__clkbuf_4 T17Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7685));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R0_INV_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7721));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R1_INV_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R2_INV_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R2_INV_1 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7757));
  sky130_fd_sc_hd__clkbuf_4 T17Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7793));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R0_INV_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7829));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R1_INV_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R2_INV_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R2_INV_1 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7865));
  sky130_fd_sc_hd__clkbuf_4 T17Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7901));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R0_INV_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7937));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R1_INV_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R2_INV_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R2_INV_1 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7973));
  sky130_fd_sc_hd__clkbuf_4 T17Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8009));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R0_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8045));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R1_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R2_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R2_INV_1 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8081));
  sky130_fd_sc_hd__clkbuf_4 T17Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8117));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R0_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8153));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R1_INV_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R2_INV_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R2_INV_1 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8189));
  sky130_fd_sc_hd__clkbuf_4 T17Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8225));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R0_INV_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8261));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R1_INV_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R2_INV_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R2_INV_1 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8297));
  sky130_fd_sc_hd__clkbuf_4 T17Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8333));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R0_INV_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8369));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R1_INV_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R2_INV_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R2_INV_1 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8405));
  sky130_fd_sc_hd__clkbuf_4 T17Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8441));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R0_INV_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8477));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R1_INV_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R2_INV_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R2_INV_1 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8513));
  sky130_fd_sc_hd__clkbuf_4 T17Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8549));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R0_INV_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8585));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R1_INV_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R2_INV_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R2_INV_1 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8621));
  sky130_fd_sc_hd__clkbuf_4 T17Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B774));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R0_INV_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B810));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R1_INV_0 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R2_INV_0 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R2_INV_1 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B846));
  sky130_fd_sc_hd__clkbuf_4 T17Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8657));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R0_INV_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8693));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R1_INV_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R2_INV_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R2_INV_1 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8729));
  sky130_fd_sc_hd__clkbuf_4 T17Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8765));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R0_INV_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8801));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R1_INV_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R2_INV_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R2_INV_1 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8837));
  sky130_fd_sc_hd__clkbuf_4 T17Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8873));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R0_INV_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8909));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R1_INV_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R2_INV_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R2_INV_1 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8945));
  sky130_fd_sc_hd__clkbuf_4 T17Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8981));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R0_INV_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9017));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R1_INV_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R2_INV_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R2_INV_1 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9053));
  sky130_fd_sc_hd__clkbuf_4 T17Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9089));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R0_INV_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9125));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R1_INV_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R2_INV_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R2_INV_1 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9161));
  sky130_fd_sc_hd__clkbuf_4 T17Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9197));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R0_INV_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9233));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R1_INV_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R2_INV_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R2_INV_1 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9269));
  sky130_fd_sc_hd__clkbuf_4 T17Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9305));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R0_INV_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9341));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R1_INV_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R2_INV_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R2_INV_1 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9377));
  sky130_fd_sc_hd__clkbuf_4 T17Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9413));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R0_INV_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9449));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R1_INV_0 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R2_INV_0 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R2_INV_1 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9485));
  sky130_fd_sc_hd__clkbuf_4 T17Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9521));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R0_INV_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9557));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R1_INV_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R2_INV_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R2_INV_1 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9593));
  sky130_fd_sc_hd__clkbuf_4 T17Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9629));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R0_INV_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9665));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R1_INV_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R2_INV_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R2_INV_1 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9701));
  sky130_fd_sc_hd__clkbuf_4 T17Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B882));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R0_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B918));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R1_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R2_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R2_INV_1 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B954));
  sky130_fd_sc_hd__clkbuf_4 T17Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B990));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R0_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1026));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R1_INV_0 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R2_INV_0 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R2_INV_1 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1062));
  sky130_fd_sc_hd__clkbuf_4 T18Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B28));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R0_INV_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B63));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R1_INV_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R2_INV_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R2_INV_1 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B98));
  sky130_fd_sc_hd__clkbuf_4 T18Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1099));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R0_INV_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1135));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R1_INV_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R2_INV_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R2_INV_1 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1171));
  sky130_fd_sc_hd__clkbuf_4 T18Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1207));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R0_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1243));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R1_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R2_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R2_INV_1 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1279));
  sky130_fd_sc_hd__clkbuf_4 T18Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1315));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R0_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1351));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R1_INV_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R2_INV_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R2_INV_1 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1387));
  sky130_fd_sc_hd__clkbuf_4 T18Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1423));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R0_INV_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1459));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R1_INV_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R2_INV_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R2_INV_1 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1495));
  sky130_fd_sc_hd__clkbuf_4 T18Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1531));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R0_INV_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1566));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R1_INV_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R2_INV_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R2_INV_1 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1602));
  sky130_fd_sc_hd__clkbuf_4 T18Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1638));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R0_INV_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1674));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R1_INV_0 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R2_INV_0 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R2_INV_1 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1710));
  sky130_fd_sc_hd__clkbuf_4 T18Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1746));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R0_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1782));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R1_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R2_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R2_INV_1 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1818));
  sky130_fd_sc_hd__clkbuf_4 T18Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1854));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R0_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1890));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R1_INV_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R2_INV_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R2_INV_1 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1926));
  sky130_fd_sc_hd__clkbuf_4 T18Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1962));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R0_INV_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1998));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R1_INV_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R2_INV_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R2_INV_1 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2034));
  sky130_fd_sc_hd__clkbuf_4 T18Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2070));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R0_INV_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2106));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R1_INV_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R2_INV_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R2_INV_1 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2142));
  sky130_fd_sc_hd__clkbuf_4 T18Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B133));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R0_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B168));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R1_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R2_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R2_INV_1 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B203));
  sky130_fd_sc_hd__clkbuf_4 T18Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2178));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R0_INV_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2214));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R1_INV_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R2_INV_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R2_INV_1 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2250));
  sky130_fd_sc_hd__clkbuf_4 T18Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2286));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R0_INV_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2322));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R1_INV_0 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R2_INV_0 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R2_INV_1 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2358));
  sky130_fd_sc_hd__clkbuf_4 T18Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2394));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R0_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2430));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R1_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R2_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R2_INV_1 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2466));
  sky130_fd_sc_hd__clkbuf_4 T18Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2502));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R0_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2538));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R1_INV_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R2_INV_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R2_INV_1 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2574));
  sky130_fd_sc_hd__clkbuf_4 T18Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2610));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R0_INV_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2646));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R1_INV_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R2_INV_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R2_INV_1 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2682));
  sky130_fd_sc_hd__clkbuf_4 T18Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2718));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R0_INV_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2754));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R1_INV_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R2_INV_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R2_INV_1 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2790));
  sky130_fd_sc_hd__clkbuf_4 T18Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2826));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R0_INV_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2862));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R1_INV_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R2_INV_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R2_INV_1 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2898));
  sky130_fd_sc_hd__clkbuf_4 T18Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2934));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R0_INV_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2970));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R1_INV_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R2_INV_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R2_INV_1 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3006));
  sky130_fd_sc_hd__clkbuf_4 T18Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3042));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R0_INV_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3078));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R1_INV_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R2_INV_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R2_INV_1 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3114));
  sky130_fd_sc_hd__clkbuf_4 T18Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3150));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R0_INV_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3186));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R1_INV_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R2_INV_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R2_INV_1 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3222));
  sky130_fd_sc_hd__clkbuf_4 T18Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B238));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R0_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B273));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R1_INV_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R2_INV_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R2_INV_1 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B309));
  sky130_fd_sc_hd__clkbuf_4 T18Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3258));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R0_INV_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3294));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R1_INV_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R2_INV_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R2_INV_1 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3330));
  sky130_fd_sc_hd__clkbuf_4 T18Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3366));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R0_INV_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3402));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R1_INV_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R2_INV_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R2_INV_1 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3438));
  sky130_fd_sc_hd__clkbuf_4 T18Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3474));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R0_INV_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3510));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R1_INV_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R2_INV_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R2_INV_1 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3546));
  sky130_fd_sc_hd__clkbuf_4 T18Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3582));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R0_INV_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3618));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R1_INV_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R2_INV_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R2_INV_1 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3654));
  sky130_fd_sc_hd__clkbuf_4 T18Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3690));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R0_INV_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3726));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R1_INV_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R2_INV_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R2_INV_1 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3762));
  sky130_fd_sc_hd__clkbuf_4 T18Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3798));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R0_INV_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3834));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R1_INV_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R2_INV_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R2_INV_1 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3870));
  sky130_fd_sc_hd__clkbuf_4 T18Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3906));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R0_INV_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3942));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R1_INV_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R2_INV_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R2_INV_1 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3978));
  sky130_fd_sc_hd__clkbuf_4 T18Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4014));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R0_INV_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4050));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R1_INV_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R2_INV_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R2_INV_1 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4086));
  sky130_fd_sc_hd__clkbuf_4 T18Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4122));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R0_INV_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4158));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R1_INV_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R2_INV_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R2_INV_1 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4194));
  sky130_fd_sc_hd__clkbuf_4 T18Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4230));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R0_INV_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4266));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R1_INV_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R2_INV_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R2_INV_1 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4302));
  sky130_fd_sc_hd__clkbuf_4 T18Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B344));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R0_INV_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B379));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R1_INV_0 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R2_INV_0 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R2_INV_1 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B415));
  sky130_fd_sc_hd__clkbuf_4 T18Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4338));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R0_INV_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4374));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R1_INV_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R2_INV_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R2_INV_1 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4410));
  sky130_fd_sc_hd__clkbuf_4 T18Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4446));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R0_INV_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4482));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R1_INV_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R2_INV_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R2_INV_1 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4518));
  sky130_fd_sc_hd__clkbuf_4 T18Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4554));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R0_INV_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4590));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R1_INV_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R2_INV_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R2_INV_1 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4626));
  sky130_fd_sc_hd__clkbuf_4 T18Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4662));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R0_INV_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4698));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R1_INV_0 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R2_INV_0 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R2_INV_1 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4734));
  sky130_fd_sc_hd__clkbuf_4 T18Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4770));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R0_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4806));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R1_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R2_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R2_INV_1 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4842));
  sky130_fd_sc_hd__clkbuf_4 T18Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4878));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R0_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4914));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R1_INV_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R2_INV_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R2_INV_1 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4950));
  sky130_fd_sc_hd__clkbuf_4 T18Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4986));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R0_INV_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5022));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R1_INV_0 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R2_INV_0 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R2_INV_1 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5058));
  sky130_fd_sc_hd__clkbuf_4 T18Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5094));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R0_INV_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5130));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R1_INV_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R2_INV_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R2_INV_1 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5166));
  sky130_fd_sc_hd__clkbuf_4 T18Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5202));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R0_INV_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5238));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R1_INV_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R2_INV_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R2_INV_1 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5274));
  sky130_fd_sc_hd__clkbuf_4 T18Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5310));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R0_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5346));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R1_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R2_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R2_INV_1 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5382));
  sky130_fd_sc_hd__clkbuf_4 T18Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B451));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R0_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B487));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R1_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R2_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R2_INV_1 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B523));
  sky130_fd_sc_hd__clkbuf_4 T18Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5418));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R0_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5454));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R1_INV_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R2_INV_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R2_INV_1 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5490));
  sky130_fd_sc_hd__clkbuf_4 T18Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5526));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R0_INV_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5562));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R1_INV_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R2_INV_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R2_INV_1 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5598));
  sky130_fd_sc_hd__clkbuf_4 T18Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5634));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R0_INV_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5670));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R1_INV_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R2_INV_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R2_INV_1 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5706));
  sky130_fd_sc_hd__clkbuf_4 T18Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5742));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R0_INV_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5778));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R1_INV_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R2_INV_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R2_INV_1 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5814));
  sky130_fd_sc_hd__clkbuf_4 T18Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5850));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R0_INV_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5886));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R1_INV_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R2_INV_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R2_INV_1 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5922));
  sky130_fd_sc_hd__clkbuf_4 T18Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5958));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R0_INV_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5994));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R1_INV_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R2_INV_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R2_INV_1 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6030));
  sky130_fd_sc_hd__clkbuf_4 T18Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6066));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R0_INV_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6102));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R1_INV_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R2_INV_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R2_INV_1 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6138));
  sky130_fd_sc_hd__clkbuf_4 T18Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6174));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R0_INV_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6210));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R1_INV_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R2_INV_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R2_INV_1 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6246));
  sky130_fd_sc_hd__clkbuf_4 T18Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6282));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R0_INV_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6318));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R1_INV_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R2_INV_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R2_INV_1 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6354));
  sky130_fd_sc_hd__clkbuf_4 T18Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6390));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R0_INV_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6426));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R1_INV_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R2_INV_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R2_INV_1 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6462));
  sky130_fd_sc_hd__clkbuf_4 T18Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B559));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R0_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B595));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R1_INV_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R2_INV_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R2_INV_1 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B631));
  sky130_fd_sc_hd__clkbuf_4 T18Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6498));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R0_INV_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6534));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R1_INV_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R2_INV_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R2_INV_1 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6570));
  sky130_fd_sc_hd__clkbuf_4 T18Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6606));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R0_INV_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6642));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R1_INV_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R2_INV_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R2_INV_1 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6678));
  sky130_fd_sc_hd__clkbuf_4 T18Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6714));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R0_INV_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6750));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R1_INV_0 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R2_INV_0 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R2_INV_1 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6786));
  sky130_fd_sc_hd__clkbuf_4 T18Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6822));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R0_INV_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6858));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R1_INV_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R2_INV_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R2_INV_1 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6894));
  sky130_fd_sc_hd__clkbuf_4 T18Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6930));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R0_INV_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6966));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R1_INV_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R2_INV_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R2_INV_1 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7002));
  sky130_fd_sc_hd__clkbuf_4 T18Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7038));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R0_INV_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7074));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R1_INV_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R2_INV_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R2_INV_1 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7110));
  sky130_fd_sc_hd__clkbuf_4 T18Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7146));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R0_INV_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7182));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R1_INV_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R2_INV_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R2_INV_1 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7218));
  sky130_fd_sc_hd__clkbuf_4 T18Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7254));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R0_INV_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7290));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R1_INV_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R2_INV_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R2_INV_1 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7326));
  sky130_fd_sc_hd__clkbuf_4 T18Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7362));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R0_INV_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7398));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R1_INV_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R2_INV_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R2_INV_1 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7434));
  sky130_fd_sc_hd__clkbuf_4 T18Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7470));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R0_INV_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7506));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R1_INV_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R2_INV_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R2_INV_1 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7542));
  sky130_fd_sc_hd__clkbuf_4 T18Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B667));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R0_INV_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B703));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R1_INV_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R2_INV_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R2_INV_1 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B739));
  sky130_fd_sc_hd__clkbuf_4 T18Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7578));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R0_INV_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7614));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R1_INV_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R2_INV_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R2_INV_1 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7650));
  sky130_fd_sc_hd__clkbuf_4 T18Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7686));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R0_INV_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7722));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R1_INV_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R2_INV_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R2_INV_1 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7758));
  sky130_fd_sc_hd__clkbuf_4 T18Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7794));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R0_INV_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7830));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R1_INV_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R2_INV_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R2_INV_1 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7866));
  sky130_fd_sc_hd__clkbuf_4 T18Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7902));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R0_INV_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7938));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R1_INV_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R2_INV_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R2_INV_1 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7974));
  sky130_fd_sc_hd__clkbuf_4 T18Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8010));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R0_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8046));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R1_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R2_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R2_INV_1 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8082));
  sky130_fd_sc_hd__clkbuf_4 T18Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8118));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R0_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8154));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R1_INV_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R2_INV_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R2_INV_1 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8190));
  sky130_fd_sc_hd__clkbuf_4 T18Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8226));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R0_INV_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8262));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R1_INV_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R2_INV_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R2_INV_1 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8298));
  sky130_fd_sc_hd__clkbuf_4 T18Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8334));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R0_INV_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8370));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R1_INV_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R2_INV_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R2_INV_1 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8406));
  sky130_fd_sc_hd__clkbuf_4 T18Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8442));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R0_INV_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8478));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R1_INV_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R2_INV_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R2_INV_1 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8514));
  sky130_fd_sc_hd__clkbuf_4 T18Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8550));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R0_INV_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8586));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R1_INV_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R2_INV_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R2_INV_1 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8622));
  sky130_fd_sc_hd__clkbuf_4 T18Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B775));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R0_INV_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B811));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R1_INV_0 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R2_INV_0 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R2_INV_1 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B847));
  sky130_fd_sc_hd__clkbuf_4 T18Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8658));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R0_INV_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8694));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R1_INV_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R2_INV_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R2_INV_1 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8730));
  sky130_fd_sc_hd__clkbuf_4 T18Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8766));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R0_INV_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8802));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R1_INV_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R2_INV_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R2_INV_1 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8838));
  sky130_fd_sc_hd__clkbuf_4 T18Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8874));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R0_INV_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8910));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R1_INV_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R2_INV_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R2_INV_1 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8946));
  sky130_fd_sc_hd__clkbuf_4 T18Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8982));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R0_INV_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9018));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R1_INV_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R2_INV_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R2_INV_1 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9054));
  sky130_fd_sc_hd__clkbuf_4 T18Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9090));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R0_INV_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9126));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R1_INV_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R2_INV_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R2_INV_1 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9162));
  sky130_fd_sc_hd__clkbuf_4 T18Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9198));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R0_INV_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9234));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R1_INV_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R2_INV_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R2_INV_1 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9270));
  sky130_fd_sc_hd__clkbuf_4 T18Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9306));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R0_INV_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9342));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R1_INV_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R2_INV_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R2_INV_1 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9378));
  sky130_fd_sc_hd__clkbuf_4 T18Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9414));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R0_INV_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9450));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R1_INV_0 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R2_INV_0 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R2_INV_1 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9486));
  sky130_fd_sc_hd__clkbuf_4 T18Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9522));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R0_INV_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9558));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R1_INV_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R2_INV_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R2_INV_1 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9594));
  sky130_fd_sc_hd__clkbuf_4 T18Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9630));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R0_INV_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9666));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R1_INV_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R2_INV_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R2_INV_1 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9702));
  sky130_fd_sc_hd__clkbuf_4 T18Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B883));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R0_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B919));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R1_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R2_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R2_INV_1 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B955));
  sky130_fd_sc_hd__clkbuf_4 T18Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B991));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R0_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1027));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R1_INV_0 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R2_INV_0 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R2_INV_1 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1063));
  sky130_fd_sc_hd__clkbuf_4 T19Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B29));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R0_INV_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y0__R1_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B4));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R1_INV_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R2_INV_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R2_INV_1 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B99));
  sky130_fd_sc_hd__clkbuf_4 T19Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1100));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R0_INV_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y10__R1_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B71));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R1_INV_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R2_INV_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R2_INV_1 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1172));
  sky130_fd_sc_hd__clkbuf_4 T19Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1208));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R0_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1244));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R1_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R2_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R2_INV_1 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y11__R3_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B5));
  sky130_fd_sc_hd__clkbuf_4 T19Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1316));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R0_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1352));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R1_INV_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R2_INV_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R2_INV_1 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1388));
  sky130_fd_sc_hd__clkbuf_4 T19Y13__R0_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B89));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R0_INV_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1460));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R1_INV_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R2_INV_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R2_INV_1 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1496));
  sky130_fd_sc_hd__clkbuf_4 T19Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1532));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R0_INV_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1567));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R1_INV_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R2_INV_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R2_INV_1 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1603));
  sky130_fd_sc_hd__clkbuf_4 T19Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1639));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R0_INV_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1675));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R1_INV_0 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R2_INV_0 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R2_INV_1 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1711));
  sky130_fd_sc_hd__clkbuf_4 T19Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1747));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R0_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1783));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R1_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R2_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R2_INV_1 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1819));
  sky130_fd_sc_hd__clkbuf_4 T19Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1855));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R0_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1891));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R1_INV_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R2_INV_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R2_INV_1 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1927));
  sky130_fd_sc_hd__clkbuf_4 T19Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1963));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R0_INV_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1999));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R1_INV_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R2_INV_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R2_INV_1 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2035));
  sky130_fd_sc_hd__clkbuf_4 T19Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2071));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R0_INV_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2107));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R1_INV_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R2_INV_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R2_INV_1 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2143));
  sky130_fd_sc_hd__clkbuf_4 T19Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B134));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R0_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B169));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R1_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R2_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R2_INV_1 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B204));
  sky130_fd_sc_hd__clkbuf_4 T19Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2179));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R0_INV_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2215));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R1_INV_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R2_INV_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R2_INV_1 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2251));
  sky130_fd_sc_hd__clkbuf_4 T19Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2287));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R0_INV_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2323));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R1_INV_0 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R2_INV_0 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R2_INV_1 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2359));
  sky130_fd_sc_hd__clkbuf_4 T19Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2395));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R0_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2431));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R1_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R2_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R2_INV_1 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2467));
  sky130_fd_sc_hd__clkbuf_4 T19Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2503));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R0_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2539));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R1_INV_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R2_INV_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R2_INV_1 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2575));
  sky130_fd_sc_hd__clkbuf_4 T19Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2611));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R0_INV_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2647));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R1_INV_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R2_INV_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R2_INV_1 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2683));
  sky130_fd_sc_hd__clkbuf_4 T19Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2719));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R0_INV_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2755));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R1_INV_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R2_INV_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R2_INV_1 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2791));
  sky130_fd_sc_hd__clkbuf_4 T19Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2827));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R0_INV_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2863));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R1_INV_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R2_INV_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R2_INV_1 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2899));
  sky130_fd_sc_hd__clkbuf_4 T19Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2935));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R0_INV_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2971));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R1_INV_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R2_INV_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R2_INV_1 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B3007));
  sky130_fd_sc_hd__clkbuf_4 T19Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3043));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R0_INV_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3079));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R1_INV_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R2_INV_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R2_INV_1 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3115));
  sky130_fd_sc_hd__clkbuf_4 T19Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3151));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R0_INV_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3187));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R1_INV_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R2_INV_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R2_INV_1 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3223));
  sky130_fd_sc_hd__clkbuf_4 T19Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B239));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R0_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B274));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R1_INV_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R2_INV_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R2_INV_1 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B310));
  sky130_fd_sc_hd__clkbuf_4 T19Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3259));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R0_INV_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3295));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R1_INV_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R2_INV_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R2_INV_1 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3331));
  sky130_fd_sc_hd__clkbuf_4 T19Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3367));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R0_INV_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3403));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R1_INV_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R2_INV_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R2_INV_1 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3439));
  sky130_fd_sc_hd__clkbuf_4 T19Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3475));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R0_INV_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3511));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R1_INV_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R2_INV_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R2_INV_1 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3547));
  sky130_fd_sc_hd__clkbuf_4 T19Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3583));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R0_INV_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3619));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R1_INV_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R2_INV_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R2_INV_1 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3655));
  sky130_fd_sc_hd__clkbuf_4 T19Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3691));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R0_INV_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3727));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R1_INV_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R2_INV_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R2_INV_1 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3763));
  sky130_fd_sc_hd__clkbuf_4 T19Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3799));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R0_INV_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3835));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R1_INV_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R2_INV_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R2_INV_1 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3871));
  sky130_fd_sc_hd__clkbuf_4 T19Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3907));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R0_INV_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3943));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R1_INV_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R2_INV_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R2_INV_1 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3979));
  sky130_fd_sc_hd__clkbuf_4 T19Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4015));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R0_INV_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4051));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R1_INV_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R2_INV_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R2_INV_1 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4087));
  sky130_fd_sc_hd__clkbuf_4 T19Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4123));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R0_INV_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4159));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R1_INV_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R2_INV_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R2_INV_1 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4195));
  sky130_fd_sc_hd__clkbuf_4 T19Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4231));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R0_INV_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4267));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R1_INV_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R2_INV_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R2_INV_1 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4303));
  sky130_fd_sc_hd__clkbuf_4 T19Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B345));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R0_INV_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B380));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R1_INV_0 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R2_INV_0 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R2_INV_1 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y3__R3_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B26));
  sky130_fd_sc_hd__clkbuf_4 T19Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4339));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R0_INV_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4375));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R1_INV_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R2_INV_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R2_INV_1 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4411));
  sky130_fd_sc_hd__clkbuf_4 T19Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4447));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R0_INV_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4483));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R1_INV_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R2_INV_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R2_INV_1 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4519));
  sky130_fd_sc_hd__clkbuf_4 T19Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4555));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R0_INV_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4591));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R1_INV_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R2_INV_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R2_INV_1 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4627));
  sky130_fd_sc_hd__clkbuf_4 T19Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4663));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R0_INV_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4699));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R1_INV_0 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R2_INV_0 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R2_INV_1 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4735));
  sky130_fd_sc_hd__clkbuf_4 T19Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4771));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R0_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4807));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R1_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R2_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R2_INV_1 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4843));
  sky130_fd_sc_hd__clkbuf_4 T19Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4879));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R0_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4915));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R1_INV_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R2_INV_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R2_INV_1 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4951));
  sky130_fd_sc_hd__clkbuf_4 T19Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4987));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R0_INV_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5023));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R1_INV_0 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R2_INV_0 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R2_INV_1 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5059));
  sky130_fd_sc_hd__clkbuf_4 T19Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5095));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R0_INV_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5131));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R1_INV_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R2_INV_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R2_INV_1 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5167));
  sky130_fd_sc_hd__clkbuf_4 T19Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5203));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R0_INV_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5239));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R1_INV_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R2_INV_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R2_INV_1 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5275));
  sky130_fd_sc_hd__clkbuf_4 T19Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5311));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R0_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5347));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R1_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R2_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R2_INV_1 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5383));
  sky130_fd_sc_hd__clkbuf_4 T19Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B452));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R0_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B488));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R1_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R2_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R2_INV_1 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B524));
  sky130_fd_sc_hd__clkbuf_4 T19Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5419));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R0_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5455));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R1_INV_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R2_INV_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R2_INV_1 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5491));
  sky130_fd_sc_hd__clkbuf_4 T19Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5527));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R0_INV_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5563));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R1_INV_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R2_INV_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R2_INV_1 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5599));
  sky130_fd_sc_hd__clkbuf_4 T19Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5635));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R0_INV_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5671));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R1_INV_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R2_INV_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R2_INV_1 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5707));
  sky130_fd_sc_hd__clkbuf_4 T19Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5743));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R0_INV_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5779));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R1_INV_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R2_INV_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R2_INV_1 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5815));
  sky130_fd_sc_hd__clkbuf_4 T19Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5851));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R0_INV_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5887));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R1_INV_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R2_INV_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R2_INV_1 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5923));
  sky130_fd_sc_hd__clkbuf_4 T19Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5959));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R0_INV_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5995));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R1_INV_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R2_INV_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R2_INV_1 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6031));
  sky130_fd_sc_hd__clkbuf_4 T19Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6067));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R0_INV_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6103));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R1_INV_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R2_INV_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R2_INV_1 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6139));
  sky130_fd_sc_hd__clkbuf_4 T19Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6175));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R0_INV_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6211));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R1_INV_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R2_INV_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R2_INV_1 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6247));
  sky130_fd_sc_hd__clkbuf_4 T19Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6283));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R0_INV_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6319));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R1_INV_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R2_INV_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R2_INV_1 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6355));
  sky130_fd_sc_hd__clkbuf_4 T19Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6391));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R0_INV_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6427));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R1_INV_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R2_INV_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R2_INV_1 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6463));
  sky130_fd_sc_hd__clkbuf_4 T19Y5__R0_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B35));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R0_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B596));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R1_INV_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R2_INV_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R2_INV_1 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B632));
  sky130_fd_sc_hd__clkbuf_4 T19Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6499));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R0_INV_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6535));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R1_INV_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R2_INV_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R2_INV_1 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6571));
  sky130_fd_sc_hd__clkbuf_4 T19Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6607));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R0_INV_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6643));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R1_INV_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R2_INV_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R2_INV_1 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6679));
  sky130_fd_sc_hd__clkbuf_4 T19Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6715));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R0_INV_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6751));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R1_INV_0 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R2_INV_0 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R2_INV_1 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6787));
  sky130_fd_sc_hd__clkbuf_4 T19Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6823));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R0_INV_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6859));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R1_INV_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R2_INV_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R2_INV_1 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6895));
  sky130_fd_sc_hd__clkbuf_4 T19Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6931));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R0_INV_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6967));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R1_INV_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R2_INV_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R2_INV_1 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7003));
  sky130_fd_sc_hd__clkbuf_4 T19Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7039));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R0_INV_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7075));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R1_INV_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R2_INV_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R2_INV_1 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7111));
  sky130_fd_sc_hd__clkbuf_4 T19Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7147));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R0_INV_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7183));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R1_INV_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R2_INV_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R2_INV_1 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7219));
  sky130_fd_sc_hd__clkbuf_4 T19Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7255));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R0_INV_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7291));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R1_INV_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R2_INV_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R2_INV_1 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7327));
  sky130_fd_sc_hd__clkbuf_4 T19Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7363));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R0_INV_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7399));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R1_INV_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R2_INV_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R2_INV_1 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7435));
  sky130_fd_sc_hd__clkbuf_4 T19Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7471));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R0_INV_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7507));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R1_INV_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R2_INV_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R2_INV_1 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7543));
  sky130_fd_sc_hd__clkbuf_4 T19Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B668));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R0_INV_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y6__R1_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B44));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R1_INV_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R2_INV_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R2_INV_1 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B740));
  sky130_fd_sc_hd__clkbuf_4 T19Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7579));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R0_INV_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7615));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R1_INV_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R2_INV_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R2_INV_1 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7651));
  sky130_fd_sc_hd__clkbuf_4 T19Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7687));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R0_INV_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7723));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R1_INV_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R2_INV_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R2_INV_1 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7759));
  sky130_fd_sc_hd__clkbuf_4 T19Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7795));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R0_INV_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7831));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R1_INV_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R2_INV_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R2_INV_1 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7867));
  sky130_fd_sc_hd__clkbuf_4 T19Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7903));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R0_INV_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7939));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R1_INV_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R2_INV_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R2_INV_1 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7975));
  sky130_fd_sc_hd__clkbuf_4 T19Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8011));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R0_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8047));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R1_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R2_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R2_INV_1 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8083));
  sky130_fd_sc_hd__clkbuf_4 T19Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8119));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R0_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8155));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R1_INV_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R2_INV_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R2_INV_1 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8191));
  sky130_fd_sc_hd__clkbuf_4 T19Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8227));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R0_INV_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8263));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R1_INV_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R2_INV_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R2_INV_1 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8299));
  sky130_fd_sc_hd__clkbuf_4 T19Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8335));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R0_INV_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8371));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R1_INV_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R2_INV_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R2_INV_1 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8407));
  sky130_fd_sc_hd__clkbuf_4 T19Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8443));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R0_INV_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8479));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R1_INV_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R2_INV_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R2_INV_1 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8515));
  sky130_fd_sc_hd__clkbuf_4 T19Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8551));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R0_INV_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8587));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R1_INV_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R2_INV_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R2_INV_1 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8623));
  sky130_fd_sc_hd__clkbuf_4 T19Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B776));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R0_INV_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B812));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R1_INV_0 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R2_INV_0 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R2_INV_1 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y7__R3_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B53));
  sky130_fd_sc_hd__clkbuf_4 T19Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8659));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R0_INV_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8695));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R1_INV_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R2_INV_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R2_INV_1 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8731));
  sky130_fd_sc_hd__clkbuf_4 T19Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8767));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R0_INV_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8803));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R1_INV_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R2_INV_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R2_INV_1 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8839));
  sky130_fd_sc_hd__clkbuf_4 T19Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8875));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R0_INV_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8911));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R1_INV_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R2_INV_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R2_INV_1 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8947));
  sky130_fd_sc_hd__clkbuf_4 T19Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8983));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R0_INV_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9019));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R1_INV_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R2_INV_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R2_INV_1 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9055));
  sky130_fd_sc_hd__clkbuf_4 T19Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9091));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R0_INV_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9127));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R1_INV_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R2_INV_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R2_INV_1 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9163));
  sky130_fd_sc_hd__clkbuf_4 T19Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9199));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R0_INV_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9235));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R1_INV_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R2_INV_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R2_INV_1 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9271));
  sky130_fd_sc_hd__clkbuf_4 T19Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9307));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R0_INV_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9343));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R1_INV_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R2_INV_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R2_INV_1 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9379));
  sky130_fd_sc_hd__clkbuf_4 T19Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9415));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R0_INV_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9451));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R1_INV_0 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R2_INV_0 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R2_INV_1 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9487));
  sky130_fd_sc_hd__clkbuf_4 T19Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9523));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R0_INV_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9559));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R1_INV_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R2_INV_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R2_INV_1 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9595));
  sky130_fd_sc_hd__clkbuf_4 T19Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9631));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R0_INV_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9667));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R1_INV_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R2_INV_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R2_INV_1 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9703));
  sky130_fd_sc_hd__clkbuf_4 T19Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B884));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R0_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B920));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R1_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R2_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R2_INV_1 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B956));
  sky130_fd_sc_hd__clkbuf_4 T19Y9__R0_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B62));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R0_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1028));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R1_INV_0 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R2_INV_0 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R2_INV_1 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1064));
  sky130_fd_sc_hd__clkbuf_4 T1Y0__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B11));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R0_INV_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y0__R1_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B46));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R1_INV_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R2_INV_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R2_INV_1 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B81));
  sky130_fd_sc_hd__clkbuf_4 T1Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1082));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R0_INV_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y10__R1_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1118));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R1_INV_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R2_INV_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R2_INV_1 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1154));
  sky130_fd_sc_hd__clkbuf_4 T1Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1190));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R0_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1226));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R1_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R2_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R2_INV_1 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y11__R3_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1262));
  sky130_fd_sc_hd__clkbuf_4 T1Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1298));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R0_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1334));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R1_INV_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R2_INV_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R2_INV_1 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1370));
  sky130_fd_sc_hd__clkbuf_4 T1Y13__R0_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1406));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R0_INV_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1442));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R1_INV_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R2_INV_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R2_INV_1 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1478));
  sky130_fd_sc_hd__clkbuf_4 T1Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1514));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R0_INV_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y14__R1_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1549));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R1_INV_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R2_INV_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R2_INV_1 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1585));
  sky130_fd_sc_hd__clkbuf_4 T1Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1621));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R0_INV_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1657));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R1_INV_0 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R2_INV_0 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R2_INV_1 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y15__R3_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1693));
  sky130_fd_sc_hd__clkbuf_4 T1Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1729));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R0_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1765));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R1_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R2_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R2_INV_1 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1801));
  sky130_fd_sc_hd__clkbuf_4 T1Y17__R0_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1837));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R0_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1873));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R1_INV_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R2_INV_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R2_INV_1 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1909));
  sky130_fd_sc_hd__clkbuf_4 T1Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1945));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R0_INV_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y18__R1_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1981));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R1_INV_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R2_INV_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R2_INV_1 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2017));
  sky130_fd_sc_hd__clkbuf_4 T1Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2053));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R0_INV_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2089));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R1_INV_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R2_INV_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R2_INV_1 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y19__R3_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2125));
  sky130_fd_sc_hd__clkbuf_4 T1Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B116));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R0_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B151));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R1_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R2_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R2_INV_1 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B186));
  sky130_fd_sc_hd__clkbuf_4 T1Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2161));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R0_INV_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2197));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R1_INV_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R2_INV_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R2_INV_1 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2233));
  sky130_fd_sc_hd__clkbuf_4 T1Y21__R0_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2269));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R0_INV_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2305));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R1_INV_0 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R2_INV_0 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R2_INV_1 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2341));
  sky130_fd_sc_hd__clkbuf_4 T1Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2377));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R0_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y22__R1_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2413));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R1_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R2_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R2_INV_1 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2449));
  sky130_fd_sc_hd__clkbuf_4 T1Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2485));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R0_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2521));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R1_INV_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R2_INV_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R2_INV_1 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y23__R3_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2557));
  sky130_fd_sc_hd__clkbuf_4 T1Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2593));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R0_INV_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2629));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R1_INV_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R2_INV_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R2_INV_1 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2665));
  sky130_fd_sc_hd__clkbuf_4 T1Y25__R0_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2701));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R0_INV_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2737));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R1_INV_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R2_INV_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R2_INV_1 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2773));
  sky130_fd_sc_hd__clkbuf_4 T1Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2809));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R0_INV_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y26__R1_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2845));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R1_INV_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R2_INV_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R2_INV_1 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2881));
  sky130_fd_sc_hd__clkbuf_4 T1Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2917));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R0_INV_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2953));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R1_INV_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R2_INV_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R2_INV_1 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y27__R3_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2989));
  sky130_fd_sc_hd__clkbuf_4 T1Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3025));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R0_INV_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3061));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R1_INV_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R2_INV_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R2_INV_1 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3097));
  sky130_fd_sc_hd__clkbuf_4 T1Y29__R0_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3133));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R0_INV_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3169));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R1_INV_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R2_INV_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R2_INV_1 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3205));
  sky130_fd_sc_hd__clkbuf_4 T1Y2__R0_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B221));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R0_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y2__R1_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B1));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R1_INV_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R2_INV_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R2_INV_1 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B292));
  sky130_fd_sc_hd__clkbuf_4 T1Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3241));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R0_INV_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y30__R1_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3277));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R1_INV_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R2_INV_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R2_INV_1 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3313));
  sky130_fd_sc_hd__clkbuf_4 T1Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3349));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R0_INV_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3385));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R1_INV_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R2_INV_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R2_INV_1 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y31__R3_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3421));
  sky130_fd_sc_hd__clkbuf_4 T1Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3457));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R0_INV_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3493));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R1_INV_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R2_INV_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R2_INV_1 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3529));
  sky130_fd_sc_hd__clkbuf_4 T1Y33__R0_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3565));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R0_INV_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3601));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R1_INV_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R2_INV_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R2_INV_1 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3637));
  sky130_fd_sc_hd__clkbuf_4 T1Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3673));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R0_INV_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y34__R1_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3709));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R1_INV_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R2_INV_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R2_INV_1 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3745));
  sky130_fd_sc_hd__clkbuf_4 T1Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3781));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R0_INV_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3817));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R1_INV_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R2_INV_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R2_INV_1 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y35__R3_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3853));
  sky130_fd_sc_hd__clkbuf_4 T1Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3889));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R0_INV_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3925));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R1_INV_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R2_INV_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R2_INV_1 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3961));
  sky130_fd_sc_hd__clkbuf_4 T1Y37__R0_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3997));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R0_INV_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4033));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R1_INV_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R2_INV_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R2_INV_1 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4069));
  sky130_fd_sc_hd__clkbuf_4 T1Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4105));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R0_INV_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y38__R1_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4141));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R1_INV_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R2_INV_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R2_INV_1 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4177));
  sky130_fd_sc_hd__clkbuf_4 T1Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4213));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R0_INV_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4249));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R1_INV_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R2_INV_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R2_INV_1 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y39__R3_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4285));
  sky130_fd_sc_hd__clkbuf_4 T1Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B327));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R0_INV_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B362));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R1_INV_0 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R2_INV_0 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R2_INV_1 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y3__R3_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B398));
  sky130_fd_sc_hd__clkbuf_4 T1Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4321));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R0_INV_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4357));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R1_INV_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R2_INV_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R2_INV_1 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4393));
  sky130_fd_sc_hd__clkbuf_4 T1Y41__R0_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4429));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R0_INV_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4465));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R1_INV_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R2_INV_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R2_INV_1 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4501));
  sky130_fd_sc_hd__clkbuf_4 T1Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4537));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R0_INV_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y42__R1_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4573));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R1_INV_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R2_INV_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R2_INV_1 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4609));
  sky130_fd_sc_hd__clkbuf_4 T1Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4645));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R0_INV_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4681));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R1_INV_0 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R2_INV_0 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R2_INV_1 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y43__R3_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4717));
  sky130_fd_sc_hd__clkbuf_4 T1Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4753));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R0_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4789));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R1_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R2_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R2_INV_1 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4825));
  sky130_fd_sc_hd__clkbuf_4 T1Y45__R0_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4861));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R0_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4897));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R1_INV_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R2_INV_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R2_INV_1 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4933));
  sky130_fd_sc_hd__clkbuf_4 T1Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4969));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R0_INV_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y46__R1_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5005));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R1_INV_0 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R2_INV_0 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R2_INV_1 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5041));
  sky130_fd_sc_hd__clkbuf_4 T1Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5077));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R0_INV_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5113));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R1_INV_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R2_INV_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R2_INV_1 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y47__R3_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5149));
  sky130_fd_sc_hd__clkbuf_4 T1Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5185));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R0_INV_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5221));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R1_INV_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R2_INV_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R2_INV_1 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5257));
  sky130_fd_sc_hd__clkbuf_4 T1Y49__R0_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5293));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R0_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5329));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R1_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R2_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R2_INV_1 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5365));
  sky130_fd_sc_hd__clkbuf_4 T1Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B434));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R0_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B470));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R1_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R2_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R2_INV_1 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B506));
  sky130_fd_sc_hd__clkbuf_4 T1Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5401));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R0_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y50__R1_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5437));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R1_INV_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R2_INV_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R2_INV_1 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5473));
  sky130_fd_sc_hd__clkbuf_4 T1Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5509));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R0_INV_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5545));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R1_INV_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R2_INV_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R2_INV_1 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y51__R3_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5581));
  sky130_fd_sc_hd__clkbuf_4 T1Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5617));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R0_INV_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5653));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R1_INV_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R2_INV_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R2_INV_1 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5689));
  sky130_fd_sc_hd__clkbuf_4 T1Y53__R0_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5725));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R0_INV_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5761));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R1_INV_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R2_INV_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R2_INV_1 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5797));
  sky130_fd_sc_hd__clkbuf_4 T1Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5833));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R0_INV_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y54__R1_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5869));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R1_INV_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R2_INV_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R2_INV_1 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5905));
  sky130_fd_sc_hd__clkbuf_4 T1Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5941));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R0_INV_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5977));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R1_INV_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R2_INV_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R2_INV_1 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y55__R3_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6013));
  sky130_fd_sc_hd__clkbuf_4 T1Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6049));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R0_INV_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6085));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R1_INV_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R2_INV_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R2_INV_1 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6121));
  sky130_fd_sc_hd__clkbuf_4 T1Y57__R0_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6157));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R0_INV_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6193));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R1_INV_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R2_INV_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R2_INV_1 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6229));
  sky130_fd_sc_hd__clkbuf_4 T1Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6265));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R0_INV_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y58__R1_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6301));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R1_INV_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R2_INV_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R2_INV_1 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6337));
  sky130_fd_sc_hd__clkbuf_4 T1Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6373));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R0_INV_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6409));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R1_INV_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R2_INV_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R2_INV_1 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y59__R3_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6445));
  sky130_fd_sc_hd__clkbuf_4 T1Y5__R0_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B542));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R0_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B578));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R1_INV_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R2_INV_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R2_INV_1 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B614));
  sky130_fd_sc_hd__clkbuf_4 T1Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6481));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R0_INV_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6517));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R1_INV_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R2_INV_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R2_INV_1 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6553));
  sky130_fd_sc_hd__clkbuf_4 T1Y61__R0_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6589));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R0_INV_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6625));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R1_INV_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R2_INV_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R2_INV_1 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6661));
  sky130_fd_sc_hd__clkbuf_4 T1Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6697));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R0_INV_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y62__R1_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6733));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R1_INV_0 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R2_INV_0 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R2_INV_1 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6769));
  sky130_fd_sc_hd__clkbuf_4 T1Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6805));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R0_INV_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6841));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R1_INV_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R2_INV_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R2_INV_1 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y63__R3_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6877));
  sky130_fd_sc_hd__clkbuf_4 T1Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6913));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R0_INV_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6949));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R1_INV_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R2_INV_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R2_INV_1 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6985));
  sky130_fd_sc_hd__clkbuf_4 T1Y65__R0_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7021));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R0_INV_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7057));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R1_INV_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R2_INV_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R2_INV_1 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7093));
  sky130_fd_sc_hd__clkbuf_4 T1Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7129));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R0_INV_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y66__R1_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7165));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R1_INV_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R2_INV_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R2_INV_1 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7201));
  sky130_fd_sc_hd__clkbuf_4 T1Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7237));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R0_INV_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7273));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R1_INV_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R2_INV_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R2_INV_1 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y67__R3_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7309));
  sky130_fd_sc_hd__clkbuf_4 T1Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7345));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R0_INV_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7381));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R1_INV_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R2_INV_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R2_INV_1 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7417));
  sky130_fd_sc_hd__clkbuf_4 T1Y69__R0_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7453));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R0_INV_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7489));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R1_INV_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R2_INV_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R2_INV_1 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7525));
  sky130_fd_sc_hd__clkbuf_4 T1Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B650));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R0_INV_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y6__R1_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B686));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R1_INV_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R2_INV_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R2_INV_1 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B722));
  sky130_fd_sc_hd__clkbuf_4 T1Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7561));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R0_INV_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y70__R1_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7597));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R1_INV_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R2_INV_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R2_INV_1 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7633));
  sky130_fd_sc_hd__clkbuf_4 T1Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7669));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R0_INV_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7705));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R1_INV_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R2_INV_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R2_INV_1 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y71__R3_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7741));
  sky130_fd_sc_hd__clkbuf_4 T1Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7777));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R0_INV_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7813));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R1_INV_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R2_INV_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R2_INV_1 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7849));
  sky130_fd_sc_hd__clkbuf_4 T1Y73__R0_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7885));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R0_INV_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7921));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R1_INV_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R2_INV_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R2_INV_1 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7957));
  sky130_fd_sc_hd__clkbuf_4 T1Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7993));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R0_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y74__R1_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8029));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R1_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R2_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R2_INV_1 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8065));
  sky130_fd_sc_hd__clkbuf_4 T1Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8101));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R0_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8137));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R1_INV_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R2_INV_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R2_INV_1 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y75__R3_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8173));
  sky130_fd_sc_hd__clkbuf_4 T1Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8209));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R0_INV_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8245));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R1_INV_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R2_INV_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R2_INV_1 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8281));
  sky130_fd_sc_hd__clkbuf_4 T1Y77__R0_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8317));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R0_INV_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8353));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R1_INV_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R2_INV_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R2_INV_1 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8389));
  sky130_fd_sc_hd__clkbuf_4 T1Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8425));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R0_INV_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y78__R1_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8461));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R1_INV_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R2_INV_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R2_INV_1 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8497));
  sky130_fd_sc_hd__clkbuf_4 T1Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8533));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R0_INV_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8569));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R1_INV_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R2_INV_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R2_INV_1 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y79__R3_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8605));
  sky130_fd_sc_hd__clkbuf_4 T1Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B758));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R0_INV_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B794));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R1_INV_0 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R2_INV_0 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R2_INV_1 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y7__R3_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B830));
  sky130_fd_sc_hd__clkbuf_4 T1Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8641));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R0_INV_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8677));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R1_INV_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R2_INV_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R2_INV_1 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8713));
  sky130_fd_sc_hd__clkbuf_4 T1Y81__R0_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8749));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R0_INV_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8785));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R1_INV_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R2_INV_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R2_INV_1 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8821));
  sky130_fd_sc_hd__clkbuf_4 T1Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8857));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R0_INV_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y82__R1_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8893));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R1_INV_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R2_INV_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R2_INV_1 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8929));
  sky130_fd_sc_hd__clkbuf_4 T1Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8965));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R0_INV_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9001));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R1_INV_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R2_INV_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R2_INV_1 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y83__R3_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9037));
  sky130_fd_sc_hd__clkbuf_4 T1Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9073));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R0_INV_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9109));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R1_INV_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R2_INV_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R2_INV_1 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9145));
  sky130_fd_sc_hd__clkbuf_4 T1Y85__R0_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9181));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R0_INV_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9217));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R1_INV_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R2_INV_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R2_INV_1 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9253));
  sky130_fd_sc_hd__clkbuf_4 T1Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9289));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R0_INV_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y86__R1_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9325));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R1_INV_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R2_INV_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R2_INV_1 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9361));
  sky130_fd_sc_hd__clkbuf_4 T1Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9397));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R0_INV_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9433));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R1_INV_0 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R2_INV_0 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R2_INV_1 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y87__R3_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9469));
  sky130_fd_sc_hd__clkbuf_4 T1Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9505));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R0_INV_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9541));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R1_INV_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R2_INV_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R2_INV_1 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9577));
  sky130_fd_sc_hd__clkbuf_4 T1Y89__R0_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9613));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R0_INV_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9649));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R1_INV_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R2_INV_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R2_INV_1 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9685));
  sky130_fd_sc_hd__clkbuf_4 T1Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B866));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R0_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B902));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R1_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R2_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R2_INV_1 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B938));
  sky130_fd_sc_hd__clkbuf_4 T1Y9__R0_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B974));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R0_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1010));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R1_INV_0 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R2_INV_0 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R2_INV_1 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1046));
  sky130_fd_sc_hd__clkbuf_4 T20Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B30));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R0_INV_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B65));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R1_INV_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R2_INV_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R2_INV_1 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B100));
  sky130_fd_sc_hd__clkbuf_4 T20Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1101));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R0_INV_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1137));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R1_INV_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R2_INV_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R2_INV_1 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1173));
  sky130_fd_sc_hd__clkbuf_4 T20Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1209));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R0_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1245));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R1_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R2_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R2_INV_1 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1281));
  sky130_fd_sc_hd__clkbuf_4 T20Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1317));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R0_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1353));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R1_INV_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R2_INV_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R2_INV_1 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1389));
  sky130_fd_sc_hd__clkbuf_4 T20Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1425));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R0_INV_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1461));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R1_INV_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R2_INV_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R2_INV_1 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1497));
  sky130_fd_sc_hd__clkbuf_4 T20Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1533));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R0_INV_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y14__R1_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B98));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R1_INV_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R2_INV_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R2_INV_1 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1604));
  sky130_fd_sc_hd__clkbuf_4 T20Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1640));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R0_INV_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1676));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R1_INV_0 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R2_INV_0 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R2_INV_1 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y15__R3_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B107));
  sky130_fd_sc_hd__clkbuf_4 T20Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1748));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R0_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1784));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R1_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R2_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R2_INV_1 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1820));
  sky130_fd_sc_hd__clkbuf_4 T20Y17__R0_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B116));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R0_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1892));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R1_INV_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R2_INV_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R2_INV_1 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1928));
  sky130_fd_sc_hd__clkbuf_4 T20Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1964));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R0_INV_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y18__R1_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B125));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R1_INV_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R2_INV_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R2_INV_1 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2036));
  sky130_fd_sc_hd__clkbuf_4 T20Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2072));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R0_INV_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2108));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R1_INV_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R2_INV_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R2_INV_1 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y19__R3_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B134));
  sky130_fd_sc_hd__clkbuf_4 T20Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B135));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R0_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B170));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R1_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R2_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R2_INV_1 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B205));
  sky130_fd_sc_hd__clkbuf_4 T20Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2180));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R0_INV_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2216));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R1_INV_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R2_INV_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R2_INV_1 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2252));
  sky130_fd_sc_hd__clkbuf_4 T20Y21__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B143));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R0_INV_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2324));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R1_INV_0 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R2_INV_0 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R2_INV_1 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2360));
  sky130_fd_sc_hd__clkbuf_4 T20Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2396));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R0_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y22__R1_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B152));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R1_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R2_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R2_INV_1 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2468));
  sky130_fd_sc_hd__clkbuf_4 T20Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2504));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R0_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2540));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R1_INV_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R2_INV_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R2_INV_1 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y23__R3_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B161));
  sky130_fd_sc_hd__clkbuf_4 T20Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2612));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R0_INV_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2648));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R1_INV_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R2_INV_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R2_INV_1 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2684));
  sky130_fd_sc_hd__clkbuf_4 T20Y25__R0_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B170));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R0_INV_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2756));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R1_INV_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R2_INV_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R2_INV_1 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2792));
  sky130_fd_sc_hd__clkbuf_4 T20Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2828));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R0_INV_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y26__R1_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B179));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R1_INV_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R2_INV_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R2_INV_1 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2900));
  sky130_fd_sc_hd__clkbuf_4 T20Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2936));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R0_INV_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2972));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R1_INV_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R2_INV_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R2_INV_1 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y27__R3_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B188));
  sky130_fd_sc_hd__clkbuf_4 T20Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3044));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R0_INV_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3080));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R1_INV_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R2_INV_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R2_INV_1 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3116));
  sky130_fd_sc_hd__clkbuf_4 T20Y29__R0_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B197));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R0_INV_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3188));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R1_INV_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R2_INV_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R2_INV_1 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3224));
  sky130_fd_sc_hd__clkbuf_4 T20Y2__R0_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B15));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R0_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B275));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R1_INV_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R2_INV_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R2_INV_1 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B311));
  sky130_fd_sc_hd__clkbuf_4 T20Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3260));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R0_INV_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y30__R1_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B206));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R1_INV_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R2_INV_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R2_INV_1 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3332));
  sky130_fd_sc_hd__clkbuf_4 T20Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3368));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R0_INV_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3404));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R1_INV_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R2_INV_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R2_INV_1 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y31__R3_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B215));
  sky130_fd_sc_hd__clkbuf_4 T20Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3476));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R0_INV_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3512));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R1_INV_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R2_INV_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R2_INV_1 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3548));
  sky130_fd_sc_hd__clkbuf_4 T20Y33__R0_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B14));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R0_INV_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3620));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R1_INV_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R2_INV_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R2_INV_1 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3656));
  sky130_fd_sc_hd__clkbuf_4 T20Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3692));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R0_INV_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y34__R1_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B233));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R1_INV_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R2_INV_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R2_INV_1 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3764));
  sky130_fd_sc_hd__clkbuf_4 T20Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3800));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R0_INV_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3836));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R1_INV_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R2_INV_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R2_INV_1 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y35__R3_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B242));
  sky130_fd_sc_hd__clkbuf_4 T20Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3908));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R0_INV_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3944));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R1_INV_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R2_INV_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R2_INV_1 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3980));
  sky130_fd_sc_hd__clkbuf_4 T20Y37__R0_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B251));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R0_INV_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4052));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R1_INV_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R2_INV_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R2_INV_1 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4088));
  sky130_fd_sc_hd__clkbuf_4 T20Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4124));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R0_INV_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y38__R1_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B260));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R1_INV_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R2_INV_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R2_INV_1 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4196));
  sky130_fd_sc_hd__clkbuf_4 T20Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4232));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R0_INV_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4268));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R1_INV_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R2_INV_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R2_INV_1 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y39__R3_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B269));
  sky130_fd_sc_hd__clkbuf_4 T20Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B346));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R0_INV_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B381));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R1_INV_0 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R2_INV_0 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R2_INV_1 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B417));
  sky130_fd_sc_hd__clkbuf_4 T20Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4340));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R0_INV_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4376));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R1_INV_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R2_INV_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R2_INV_1 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4412));
  sky130_fd_sc_hd__clkbuf_4 T20Y41__R0_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B278));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R0_INV_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4484));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R1_INV_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R2_INV_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R2_INV_1 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4520));
  sky130_fd_sc_hd__clkbuf_4 T20Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4556));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R0_INV_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y42__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B287));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R1_INV_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R2_INV_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R2_INV_1 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4628));
  sky130_fd_sc_hd__clkbuf_4 T20Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4664));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R0_INV_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4700));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R1_INV_0 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R2_INV_0 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R2_INV_1 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y43__R3_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B296));
  sky130_fd_sc_hd__clkbuf_4 T20Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4772));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R0_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4808));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R1_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R2_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R2_INV_1 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4844));
  sky130_fd_sc_hd__clkbuf_4 T20Y45__R0_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B305));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R0_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4916));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R1_INV_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R2_INV_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R2_INV_1 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4952));
  sky130_fd_sc_hd__clkbuf_4 T20Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4988));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R0_INV_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y46__R1_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B314));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R1_INV_0 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R2_INV_0 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R2_INV_1 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5060));
  sky130_fd_sc_hd__clkbuf_4 T20Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5096));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R0_INV_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5132));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R1_INV_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R2_INV_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R2_INV_1 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y47__R3_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B323));
  sky130_fd_sc_hd__clkbuf_4 T20Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5204));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R0_INV_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5240));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R1_INV_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R2_INV_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R2_INV_1 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5276));
  sky130_fd_sc_hd__clkbuf_4 T20Y49__R0_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B332));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R0_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5348));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R1_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R2_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R2_INV_1 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5384));
  sky130_fd_sc_hd__clkbuf_4 T20Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B453));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R0_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B489));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R1_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R2_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R2_INV_1 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B525));
  sky130_fd_sc_hd__clkbuf_4 T20Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5420));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R0_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y50__R1_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B341));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R1_INV_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R2_INV_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R2_INV_1 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5492));
  sky130_fd_sc_hd__clkbuf_4 T20Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5528));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R0_INV_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5564));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R1_INV_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R2_INV_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R2_INV_1 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y51__R3_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B350));
  sky130_fd_sc_hd__clkbuf_4 T20Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5636));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R0_INV_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5672));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R1_INV_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R2_INV_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R2_INV_1 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5708));
  sky130_fd_sc_hd__clkbuf_4 T20Y53__R0_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B359));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R0_INV_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5780));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R1_INV_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R2_INV_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R2_INV_1 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5816));
  sky130_fd_sc_hd__clkbuf_4 T20Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5852));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R0_INV_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y54__R1_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B23));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R1_INV_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R2_INV_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R2_INV_1 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5924));
  sky130_fd_sc_hd__clkbuf_4 T20Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5960));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R0_INV_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5996));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R1_INV_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R2_INV_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R2_INV_1 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y55__R3_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B377));
  sky130_fd_sc_hd__clkbuf_4 T20Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6068));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R0_INV_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6104));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R1_INV_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R2_INV_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R2_INV_1 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6140));
  sky130_fd_sc_hd__clkbuf_4 T20Y57__R0_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B386));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R0_INV_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6212));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R1_INV_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R2_INV_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R2_INV_1 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6248));
  sky130_fd_sc_hd__clkbuf_4 T20Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6284));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R0_INV_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y58__R1_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B395));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R1_INV_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R2_INV_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R2_INV_1 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6356));
  sky130_fd_sc_hd__clkbuf_4 T20Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6392));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R0_INV_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6428));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R1_INV_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R2_INV_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R2_INV_1 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y59__R3_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B404));
  sky130_fd_sc_hd__clkbuf_4 T20Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B561));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R0_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B597));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R1_INV_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R2_INV_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R2_INV_1 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B633));
  sky130_fd_sc_hd__clkbuf_4 T20Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6500));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R0_INV_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6536));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R1_INV_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R2_INV_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R2_INV_1 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6572));
  sky130_fd_sc_hd__clkbuf_4 T20Y61__R0_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B413));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R0_INV_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6644));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R1_INV_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R2_INV_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R2_INV_1 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6680));
  sky130_fd_sc_hd__clkbuf_4 T20Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6716));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R0_INV_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y62__R1_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B422));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R1_INV_0 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R2_INV_0 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R2_INV_1 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6788));
  sky130_fd_sc_hd__clkbuf_4 T20Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6824));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R0_INV_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6860));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R1_INV_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R2_INV_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R2_INV_1 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y63__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B431));
  sky130_fd_sc_hd__clkbuf_4 T20Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6932));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R0_INV_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6968));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R1_INV_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R2_INV_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R2_INV_1 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7004));
  sky130_fd_sc_hd__clkbuf_4 T20Y65__R0_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B440));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R0_INV_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7076));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R1_INV_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R2_INV_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R2_INV_1 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7112));
  sky130_fd_sc_hd__clkbuf_4 T20Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7148));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R0_INV_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y66__R1_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B449));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R1_INV_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R2_INV_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R2_INV_1 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7220));
  sky130_fd_sc_hd__clkbuf_4 T20Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7256));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R0_INV_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7292));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R1_INV_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R2_INV_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R2_INV_1 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y67__R3_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B458));
  sky130_fd_sc_hd__clkbuf_4 T20Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7364));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R0_INV_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7400));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R1_INV_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R2_INV_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R2_INV_1 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7436));
  sky130_fd_sc_hd__clkbuf_4 T20Y69__R0_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B467));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R0_INV_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7508));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R1_INV_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R2_INV_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R2_INV_1 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7544));
  sky130_fd_sc_hd__clkbuf_4 T20Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B669));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R0_INV_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B705));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R1_INV_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R2_INV_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R2_INV_1 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B741));
  sky130_fd_sc_hd__clkbuf_4 T20Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7580));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R0_INV_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y70__R1_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B476));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R1_INV_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R2_INV_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R2_INV_1 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7652));
  sky130_fd_sc_hd__clkbuf_4 T20Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7688));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R0_INV_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7724));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R1_INV_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R2_INV_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R2_INV_1 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y71__R3_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B485));
  sky130_fd_sc_hd__clkbuf_4 T20Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7796));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R0_INV_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7832));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R1_INV_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R2_INV_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R2_INV_1 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7868));
  sky130_fd_sc_hd__clkbuf_4 T20Y73__R0_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B494));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R0_INV_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7940));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R1_INV_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R2_INV_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R2_INV_1 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7976));
  sky130_fd_sc_hd__clkbuf_4 T20Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8012));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R0_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y74__R1_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B503));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R1_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R2_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R2_INV_1 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8084));
  sky130_fd_sc_hd__clkbuf_4 T20Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8120));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R0_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8156));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R1_INV_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R2_INV_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R2_INV_1 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y75__R3_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B32));
  sky130_fd_sc_hd__clkbuf_4 T20Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8228));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R0_INV_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8264));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R1_INV_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R2_INV_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R2_INV_1 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8300));
  sky130_fd_sc_hd__clkbuf_4 T20Y77__R0_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B521));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R0_INV_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8372));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R1_INV_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R2_INV_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R2_INV_1 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8408));
  sky130_fd_sc_hd__clkbuf_4 T20Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8444));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R0_INV_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y78__R1_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B530));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R1_INV_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R2_INV_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R2_INV_1 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8516));
  sky130_fd_sc_hd__clkbuf_4 T20Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8552));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R0_INV_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8588));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R1_INV_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R2_INV_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R2_INV_1 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y79__R3_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B539));
  sky130_fd_sc_hd__clkbuf_4 T20Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B777));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R0_INV_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B813));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R1_INV_0 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R2_INV_0 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R2_INV_1 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B849));
  sky130_fd_sc_hd__clkbuf_4 T20Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8660));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R0_INV_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8696));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R1_INV_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R2_INV_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R2_INV_1 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8732));
  sky130_fd_sc_hd__clkbuf_4 T20Y81__R0_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B548));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R0_INV_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8804));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R1_INV_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R2_INV_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R2_INV_1 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8840));
  sky130_fd_sc_hd__clkbuf_4 T20Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8876));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R0_INV_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y82__R1_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B557));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R1_INV_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R2_INV_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R2_INV_1 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8948));
  sky130_fd_sc_hd__clkbuf_4 T20Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8984));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R0_INV_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9020));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R1_INV_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R2_INV_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R2_INV_1 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y83__R3_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B566));
  sky130_fd_sc_hd__clkbuf_4 T20Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9092));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R0_INV_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9128));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R1_INV_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R2_INV_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R2_INV_1 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9164));
  sky130_fd_sc_hd__clkbuf_4 T20Y85__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B575));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R0_INV_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9236));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R1_INV_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R2_INV_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R2_INV_1 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9272));
  sky130_fd_sc_hd__clkbuf_4 T20Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9308));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R0_INV_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y86__R1_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B584));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R1_INV_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R2_INV_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R2_INV_1 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9380));
  sky130_fd_sc_hd__clkbuf_4 T20Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9416));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R0_INV_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9452));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R1_INV_0 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R2_INV_0 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R2_INV_1 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y87__R3_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B593));
  sky130_fd_sc_hd__clkbuf_4 T20Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9524));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R0_INV_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9560));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R1_INV_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R2_INV_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R2_INV_1 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9596));
  sky130_fd_sc_hd__clkbuf_4 T20Y89__R0_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B602));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R0_INV_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9668));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R1_INV_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R2_INV_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R2_INV_1 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9704));
  sky130_fd_sc_hd__clkbuf_4 T20Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B885));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R0_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B921));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R1_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R2_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R2_INV_1 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B957));
  sky130_fd_sc_hd__clkbuf_4 T20Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B993));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R0_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1029));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R1_INV_0 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R2_INV_0 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R2_INV_1 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1065));
  sky130_fd_sc_hd__clkbuf_4 T21Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B31));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R0_INV_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B66));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R1_INV_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R2_INV_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R2_INV_1 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B101));
  sky130_fd_sc_hd__clkbuf_4 T21Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1102));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R0_INV_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1138));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R1_INV_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R2_INV_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R2_INV_1 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1174));
  sky130_fd_sc_hd__clkbuf_4 T21Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1210));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R0_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1246));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R1_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R2_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R2_INV_1 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1282));
  sky130_fd_sc_hd__clkbuf_4 T21Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1318));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R0_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1354));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R1_INV_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R2_INV_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R2_INV_1 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1390));
  sky130_fd_sc_hd__clkbuf_4 T21Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1426));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R0_INV_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1462));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R1_INV_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R2_INV_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R2_INV_1 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1498));
  sky130_fd_sc_hd__clkbuf_4 T21Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1534));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R0_INV_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1569));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R1_INV_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R2_INV_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R2_INV_1 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1605));
  sky130_fd_sc_hd__clkbuf_4 T21Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1641));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R0_INV_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1677));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R1_INV_0 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R2_INV_0 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R2_INV_1 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1713));
  sky130_fd_sc_hd__clkbuf_4 T21Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1749));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R0_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1785));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R1_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R2_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R2_INV_1 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1821));
  sky130_fd_sc_hd__clkbuf_4 T21Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1857));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R0_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1893));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R1_INV_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R2_INV_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R2_INV_1 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1929));
  sky130_fd_sc_hd__clkbuf_4 T21Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1965));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R0_INV_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2001));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R1_INV_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R2_INV_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R2_INV_1 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2037));
  sky130_fd_sc_hd__clkbuf_4 T21Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2073));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R0_INV_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2109));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R1_INV_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R2_INV_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R2_INV_1 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2145));
  sky130_fd_sc_hd__clkbuf_4 T21Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B136));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R0_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B171));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R1_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R2_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R2_INV_1 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B206));
  sky130_fd_sc_hd__clkbuf_4 T21Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2181));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R0_INV_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2217));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R1_INV_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R2_INV_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R2_INV_1 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2253));
  sky130_fd_sc_hd__clkbuf_4 T21Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2289));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R0_INV_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2325));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R1_INV_0 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R2_INV_0 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R2_INV_1 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2361));
  sky130_fd_sc_hd__clkbuf_4 T21Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2397));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R0_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2433));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R1_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R2_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R2_INV_1 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2469));
  sky130_fd_sc_hd__clkbuf_4 T21Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2505));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R0_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2541));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R1_INV_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R2_INV_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R2_INV_1 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2577));
  sky130_fd_sc_hd__clkbuf_4 T21Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2613));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R0_INV_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2649));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R1_INV_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R2_INV_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R2_INV_1 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2685));
  sky130_fd_sc_hd__clkbuf_4 T21Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2721));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R0_INV_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2757));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R1_INV_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R2_INV_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R2_INV_1 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2793));
  sky130_fd_sc_hd__clkbuf_4 T21Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2829));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R0_INV_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2865));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R1_INV_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R2_INV_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R2_INV_1 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2901));
  sky130_fd_sc_hd__clkbuf_4 T21Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2937));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R0_INV_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2973));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R1_INV_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R2_INV_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R2_INV_1 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3009));
  sky130_fd_sc_hd__clkbuf_4 T21Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3045));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R0_INV_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3081));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R1_INV_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R2_INV_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R2_INV_1 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3117));
  sky130_fd_sc_hd__clkbuf_4 T21Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3153));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R0_INV_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3189));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R1_INV_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R2_INV_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R2_INV_1 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3225));
  sky130_fd_sc_hd__clkbuf_4 T21Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B241));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R0_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B276));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R1_INV_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R2_INV_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R2_INV_1 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B312));
  sky130_fd_sc_hd__clkbuf_4 T21Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3261));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R0_INV_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3297));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R1_INV_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R2_INV_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R2_INV_1 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3333));
  sky130_fd_sc_hd__clkbuf_4 T21Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3369));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R0_INV_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3405));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R1_INV_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R2_INV_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R2_INV_1 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3441));
  sky130_fd_sc_hd__clkbuf_4 T21Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3477));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R0_INV_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3513));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R1_INV_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R2_INV_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R2_INV_1 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3549));
  sky130_fd_sc_hd__clkbuf_4 T21Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3585));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R0_INV_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3621));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R1_INV_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R2_INV_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R2_INV_1 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3657));
  sky130_fd_sc_hd__clkbuf_4 T21Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3693));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R0_INV_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3729));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R1_INV_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R2_INV_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R2_INV_1 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3765));
  sky130_fd_sc_hd__clkbuf_4 T21Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3801));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R0_INV_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3837));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R1_INV_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R2_INV_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R2_INV_1 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3873));
  sky130_fd_sc_hd__clkbuf_4 T21Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3909));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R0_INV_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3945));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R1_INV_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R2_INV_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R2_INV_1 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3981));
  sky130_fd_sc_hd__clkbuf_4 T21Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4017));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R0_INV_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4053));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R1_INV_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R2_INV_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R2_INV_1 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4089));
  sky130_fd_sc_hd__clkbuf_4 T21Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4125));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R0_INV_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4161));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R1_INV_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R2_INV_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R2_INV_1 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4197));
  sky130_fd_sc_hd__clkbuf_4 T21Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4233));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R0_INV_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4269));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R1_INV_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R2_INV_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R2_INV_1 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4305));
  sky130_fd_sc_hd__clkbuf_4 T21Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B347));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R0_INV_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B382));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R1_INV_0 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R2_INV_0 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R2_INV_1 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B418));
  sky130_fd_sc_hd__clkbuf_4 T21Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4341));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R0_INV_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4377));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R1_INV_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R2_INV_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R2_INV_1 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4413));
  sky130_fd_sc_hd__clkbuf_4 T21Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4449));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R0_INV_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4485));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R1_INV_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R2_INV_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R2_INV_1 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4521));
  sky130_fd_sc_hd__clkbuf_4 T21Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4557));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R0_INV_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4593));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R1_INV_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R2_INV_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R2_INV_1 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4629));
  sky130_fd_sc_hd__clkbuf_4 T21Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4665));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R0_INV_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4701));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R1_INV_0 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R2_INV_0 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R2_INV_1 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4737));
  sky130_fd_sc_hd__clkbuf_4 T21Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4773));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R0_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4809));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R1_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R2_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R2_INV_1 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4845));
  sky130_fd_sc_hd__clkbuf_4 T21Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4881));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R0_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4917));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R1_INV_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R2_INV_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R2_INV_1 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4953));
  sky130_fd_sc_hd__clkbuf_4 T21Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4989));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R0_INV_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5025));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R1_INV_0 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R2_INV_0 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R2_INV_1 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5061));
  sky130_fd_sc_hd__clkbuf_4 T21Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5097));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R0_INV_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5133));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R1_INV_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R2_INV_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R2_INV_1 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5169));
  sky130_fd_sc_hd__clkbuf_4 T21Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5205));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R0_INV_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5241));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R1_INV_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R2_INV_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R2_INV_1 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5277));
  sky130_fd_sc_hd__clkbuf_4 T21Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5313));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R0_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5349));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R1_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R2_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R2_INV_1 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5385));
  sky130_fd_sc_hd__clkbuf_4 T21Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B454));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R0_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B490));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R1_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R2_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R2_INV_1 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B526));
  sky130_fd_sc_hd__clkbuf_4 T21Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5421));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R0_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5457));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R1_INV_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R2_INV_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R2_INV_1 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5493));
  sky130_fd_sc_hd__clkbuf_4 T21Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5529));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R0_INV_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5565));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R1_INV_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R2_INV_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R2_INV_1 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5601));
  sky130_fd_sc_hd__clkbuf_4 T21Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5637));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R0_INV_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5673));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R1_INV_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R2_INV_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R2_INV_1 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5709));
  sky130_fd_sc_hd__clkbuf_4 T21Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5745));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R0_INV_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5781));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R1_INV_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R2_INV_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R2_INV_1 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5817));
  sky130_fd_sc_hd__clkbuf_4 T21Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5853));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R0_INV_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5889));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R1_INV_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R2_INV_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R2_INV_1 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5925));
  sky130_fd_sc_hd__clkbuf_4 T21Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5961));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R0_INV_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5997));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R1_INV_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R2_INV_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R2_INV_1 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6033));
  sky130_fd_sc_hd__clkbuf_4 T21Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6069));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R0_INV_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6105));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R1_INV_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R2_INV_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R2_INV_1 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6141));
  sky130_fd_sc_hd__clkbuf_4 T21Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6177));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R0_INV_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6213));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R1_INV_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R2_INV_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R2_INV_1 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6249));
  sky130_fd_sc_hd__clkbuf_4 T21Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6285));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R0_INV_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6321));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R1_INV_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R2_INV_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R2_INV_1 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6357));
  sky130_fd_sc_hd__clkbuf_4 T21Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6393));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R0_INV_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6429));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R1_INV_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R2_INV_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R2_INV_1 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6465));
  sky130_fd_sc_hd__clkbuf_4 T21Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B562));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R0_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B598));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R1_INV_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R2_INV_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R2_INV_1 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B634));
  sky130_fd_sc_hd__clkbuf_4 T21Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6501));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R0_INV_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6537));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R1_INV_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R2_INV_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R2_INV_1 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6573));
  sky130_fd_sc_hd__clkbuf_4 T21Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6609));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R0_INV_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6645));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R1_INV_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R2_INV_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R2_INV_1 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6681));
  sky130_fd_sc_hd__clkbuf_4 T21Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6717));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R0_INV_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6753));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R1_INV_0 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R2_INV_0 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R2_INV_1 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6789));
  sky130_fd_sc_hd__clkbuf_4 T21Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6825));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R0_INV_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6861));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R1_INV_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R2_INV_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R2_INV_1 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6897));
  sky130_fd_sc_hd__clkbuf_4 T21Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6933));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R0_INV_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6969));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R1_INV_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R2_INV_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R2_INV_1 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7005));
  sky130_fd_sc_hd__clkbuf_4 T21Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7041));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R0_INV_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7077));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R1_INV_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R2_INV_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R2_INV_1 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7113));
  sky130_fd_sc_hd__clkbuf_4 T21Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7149));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R0_INV_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7185));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R1_INV_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R2_INV_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R2_INV_1 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7221));
  sky130_fd_sc_hd__clkbuf_4 T21Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7257));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R0_INV_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7293));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R1_INV_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R2_INV_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R2_INV_1 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7329));
  sky130_fd_sc_hd__clkbuf_4 T21Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7365));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R0_INV_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7401));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R1_INV_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R2_INV_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R2_INV_1 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7437));
  sky130_fd_sc_hd__clkbuf_4 T21Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7473));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R0_INV_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7509));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R1_INV_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R2_INV_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R2_INV_1 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7545));
  sky130_fd_sc_hd__clkbuf_4 T21Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B670));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R0_INV_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B706));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R1_INV_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R2_INV_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R2_INV_1 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B742));
  sky130_fd_sc_hd__clkbuf_4 T21Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7581));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R0_INV_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7617));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R1_INV_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R2_INV_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R2_INV_1 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7653));
  sky130_fd_sc_hd__clkbuf_4 T21Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7689));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R0_INV_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7725));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R1_INV_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R2_INV_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R2_INV_1 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7761));
  sky130_fd_sc_hd__clkbuf_4 T21Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7797));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R0_INV_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7833));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R1_INV_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R2_INV_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R2_INV_1 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7869));
  sky130_fd_sc_hd__clkbuf_4 T21Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7905));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R0_INV_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7941));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R1_INV_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R2_INV_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R2_INV_1 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7977));
  sky130_fd_sc_hd__clkbuf_4 T21Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8013));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R0_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8049));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R1_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R2_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R2_INV_1 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8085));
  sky130_fd_sc_hd__clkbuf_4 T21Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8121));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R0_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8157));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R1_INV_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R2_INV_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R2_INV_1 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8193));
  sky130_fd_sc_hd__clkbuf_4 T21Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8229));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R0_INV_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8265));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R1_INV_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R2_INV_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R2_INV_1 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8301));
  sky130_fd_sc_hd__clkbuf_4 T21Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8337));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R0_INV_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8373));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R1_INV_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R2_INV_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R2_INV_1 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8409));
  sky130_fd_sc_hd__clkbuf_4 T21Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8445));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R0_INV_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8481));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R1_INV_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R2_INV_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R2_INV_1 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8517));
  sky130_fd_sc_hd__clkbuf_4 T21Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8553));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R0_INV_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8589));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R1_INV_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R2_INV_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R2_INV_1 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8625));
  sky130_fd_sc_hd__clkbuf_4 T21Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B778));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R0_INV_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B814));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R1_INV_0 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R2_INV_0 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R2_INV_1 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B850));
  sky130_fd_sc_hd__clkbuf_4 T21Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8661));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R0_INV_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8697));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R1_INV_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R2_INV_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R2_INV_1 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8733));
  sky130_fd_sc_hd__clkbuf_4 T21Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8769));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R0_INV_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8805));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R1_INV_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R2_INV_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R2_INV_1 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8841));
  sky130_fd_sc_hd__clkbuf_4 T21Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8877));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R0_INV_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8913));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R1_INV_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R2_INV_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R2_INV_1 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8949));
  sky130_fd_sc_hd__clkbuf_4 T21Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8985));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R0_INV_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9021));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R1_INV_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R2_INV_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R2_INV_1 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9057));
  sky130_fd_sc_hd__clkbuf_4 T21Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9093));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R0_INV_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9129));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R1_INV_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R2_INV_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R2_INV_1 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9165));
  sky130_fd_sc_hd__clkbuf_4 T21Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9201));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R0_INV_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9237));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R1_INV_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R2_INV_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R2_INV_1 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9273));
  sky130_fd_sc_hd__clkbuf_4 T21Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9309));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R0_INV_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9345));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R1_INV_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R2_INV_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R2_INV_1 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9381));
  sky130_fd_sc_hd__clkbuf_4 T21Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9417));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R0_INV_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9453));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R1_INV_0 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R2_INV_0 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R2_INV_1 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9489));
  sky130_fd_sc_hd__clkbuf_4 T21Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9525));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R0_INV_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9561));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R1_INV_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R2_INV_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R2_INV_1 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9597));
  sky130_fd_sc_hd__clkbuf_4 T21Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9633));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R0_INV_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9669));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R1_INV_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R2_INV_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R2_INV_1 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9705));
  sky130_fd_sc_hd__clkbuf_4 T21Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B886));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R0_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B922));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R1_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R2_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R2_INV_1 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B958));
  sky130_fd_sc_hd__clkbuf_4 T21Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B994));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R0_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1030));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R1_INV_0 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R2_INV_0 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R2_INV_1 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1066));
  sky130_fd_sc_hd__clkbuf_4 T22Y0__R0_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B2));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R0_INV_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B67));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R1_INV_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R2_INV_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R2_INV_1 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B102));
  sky130_fd_sc_hd__clkbuf_4 T22Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1103));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R0_INV_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1139));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R1_INV_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R2_INV_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R2_INV_1 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1175));
  sky130_fd_sc_hd__clkbuf_4 T22Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1211));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R0_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1247));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R1_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R2_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R2_INV_1 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1283));
  sky130_fd_sc_hd__clkbuf_4 T22Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1319));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R0_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1355));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R1_INV_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R2_INV_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R2_INV_1 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1391));
  sky130_fd_sc_hd__clkbuf_4 T22Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1427));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R0_INV_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1463));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R1_INV_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R2_INV_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R2_INV_1 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1499));
  sky130_fd_sc_hd__clkbuf_4 T22Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1535));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R0_INV_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1570));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R1_INV_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R2_INV_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R2_INV_1 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1606));
  sky130_fd_sc_hd__clkbuf_4 T22Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1642));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R0_INV_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1678));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R1_INV_0 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R2_INV_0 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R2_INV_1 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1714));
  sky130_fd_sc_hd__clkbuf_4 T22Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1750));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R0_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1786));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R1_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R2_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R2_INV_1 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1822));
  sky130_fd_sc_hd__clkbuf_4 T22Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1858));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R0_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1894));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R1_INV_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R2_INV_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R2_INV_1 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1930));
  sky130_fd_sc_hd__clkbuf_4 T22Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1966));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R0_INV_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2002));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R1_INV_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R2_INV_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R2_INV_1 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2038));
  sky130_fd_sc_hd__clkbuf_4 T22Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2074));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R0_INV_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2110));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R1_INV_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R2_INV_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R2_INV_1 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2146));
  sky130_fd_sc_hd__clkbuf_4 T22Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B137));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R0_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B172));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R1_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R2_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R2_INV_1 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B207));
  sky130_fd_sc_hd__clkbuf_4 T22Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2182));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R0_INV_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2218));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R1_INV_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R2_INV_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R2_INV_1 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2254));
  sky130_fd_sc_hd__clkbuf_4 T22Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2290));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R0_INV_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2326));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R1_INV_0 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R2_INV_0 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R2_INV_1 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2362));
  sky130_fd_sc_hd__clkbuf_4 T22Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2398));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R0_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2434));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R1_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R2_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R2_INV_1 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2470));
  sky130_fd_sc_hd__clkbuf_4 T22Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2506));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R0_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2542));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R1_INV_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R2_INV_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R2_INV_1 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2578));
  sky130_fd_sc_hd__clkbuf_4 T22Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2614));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R0_INV_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2650));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R1_INV_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R2_INV_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R2_INV_1 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2686));
  sky130_fd_sc_hd__clkbuf_4 T22Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2722));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R0_INV_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2758));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R1_INV_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R2_INV_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R2_INV_1 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2794));
  sky130_fd_sc_hd__clkbuf_4 T22Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2830));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R0_INV_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2866));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R1_INV_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R2_INV_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R2_INV_1 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2902));
  sky130_fd_sc_hd__clkbuf_4 T22Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2938));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R0_INV_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2974));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R1_INV_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R2_INV_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R2_INV_1 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3010));
  sky130_fd_sc_hd__clkbuf_4 T22Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3046));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R0_INV_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3082));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R1_INV_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R2_INV_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R2_INV_1 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3118));
  sky130_fd_sc_hd__clkbuf_4 T22Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3154));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R0_INV_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3190));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R1_INV_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R2_INV_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R2_INV_1 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3226));
  sky130_fd_sc_hd__clkbuf_4 T22Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B242));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R0_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B277));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R1_INV_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R2_INV_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R2_INV_1 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B313));
  sky130_fd_sc_hd__clkbuf_4 T22Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3262));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R0_INV_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3298));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R1_INV_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R2_INV_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R2_INV_1 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3334));
  sky130_fd_sc_hd__clkbuf_4 T22Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3370));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R0_INV_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3406));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R1_INV_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R2_INV_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R2_INV_1 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3442));
  sky130_fd_sc_hd__clkbuf_4 T22Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3478));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R0_INV_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3514));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R1_INV_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R2_INV_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R2_INV_1 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3550));
  sky130_fd_sc_hd__clkbuf_4 T22Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3586));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R0_INV_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3622));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R1_INV_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R2_INV_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R2_INV_1 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3658));
  sky130_fd_sc_hd__clkbuf_4 T22Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3694));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R0_INV_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3730));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R1_INV_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R2_INV_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R2_INV_1 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3766));
  sky130_fd_sc_hd__clkbuf_4 T22Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3802));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R0_INV_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3838));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R1_INV_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R2_INV_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R2_INV_1 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3874));
  sky130_fd_sc_hd__clkbuf_4 T22Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3910));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R0_INV_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3946));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R1_INV_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R2_INV_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R2_INV_1 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3982));
  sky130_fd_sc_hd__clkbuf_4 T22Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4018));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R0_INV_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4054));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R1_INV_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R2_INV_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R2_INV_1 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4090));
  sky130_fd_sc_hd__clkbuf_4 T22Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4126));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R0_INV_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4162));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R1_INV_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R2_INV_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R2_INV_1 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4198));
  sky130_fd_sc_hd__clkbuf_4 T22Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4234));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R0_INV_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4270));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R1_INV_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R2_INV_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R2_INV_1 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4306));
  sky130_fd_sc_hd__clkbuf_4 T22Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B348));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R0_INV_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B383));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R1_INV_0 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R2_INV_0 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R2_INV_1 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B419));
  sky130_fd_sc_hd__clkbuf_4 T22Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4342));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R0_INV_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4378));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R1_INV_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R2_INV_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R2_INV_1 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4414));
  sky130_fd_sc_hd__clkbuf_4 T22Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4450));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R0_INV_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4486));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R1_INV_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R2_INV_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R2_INV_1 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4522));
  sky130_fd_sc_hd__clkbuf_4 T22Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4558));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R0_INV_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4594));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R1_INV_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R2_INV_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R2_INV_1 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4630));
  sky130_fd_sc_hd__clkbuf_4 T22Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4666));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R0_INV_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4702));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R1_INV_0 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R2_INV_0 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R2_INV_1 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4738));
  sky130_fd_sc_hd__clkbuf_4 T22Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4774));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R0_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4810));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R1_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R2_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R2_INV_1 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4846));
  sky130_fd_sc_hd__clkbuf_4 T22Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4882));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R0_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4918));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R1_INV_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R2_INV_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R2_INV_1 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4954));
  sky130_fd_sc_hd__clkbuf_4 T22Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4990));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R0_INV_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5026));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R1_INV_0 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R2_INV_0 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R2_INV_1 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5062));
  sky130_fd_sc_hd__clkbuf_4 T22Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5098));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R0_INV_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5134));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R1_INV_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R2_INV_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R2_INV_1 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5170));
  sky130_fd_sc_hd__clkbuf_4 T22Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5206));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R0_INV_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5242));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R1_INV_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R2_INV_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R2_INV_1 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5278));
  sky130_fd_sc_hd__clkbuf_4 T22Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5314));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R0_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5350));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R1_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R2_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R2_INV_1 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5386));
  sky130_fd_sc_hd__clkbuf_4 T22Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B455));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R0_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B491));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R1_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R2_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R2_INV_1 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B527));
  sky130_fd_sc_hd__clkbuf_4 T22Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5422));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R0_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5458));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R1_INV_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R2_INV_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R2_INV_1 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5494));
  sky130_fd_sc_hd__clkbuf_4 T22Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5530));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R0_INV_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5566));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R1_INV_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R2_INV_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R2_INV_1 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5602));
  sky130_fd_sc_hd__clkbuf_4 T22Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5638));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R0_INV_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5674));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R1_INV_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R2_INV_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R2_INV_1 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5710));
  sky130_fd_sc_hd__clkbuf_4 T22Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5746));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R0_INV_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5782));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R1_INV_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R2_INV_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R2_INV_1 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5818));
  sky130_fd_sc_hd__clkbuf_4 T22Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5854));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R0_INV_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5890));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R1_INV_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R2_INV_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R2_INV_1 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5926));
  sky130_fd_sc_hd__clkbuf_4 T22Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5962));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R0_INV_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5998));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R1_INV_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R2_INV_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R2_INV_1 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6034));
  sky130_fd_sc_hd__clkbuf_4 T22Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6070));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R0_INV_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6106));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R1_INV_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R2_INV_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R2_INV_1 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6142));
  sky130_fd_sc_hd__clkbuf_4 T22Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6178));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R0_INV_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6214));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R1_INV_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R2_INV_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R2_INV_1 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6250));
  sky130_fd_sc_hd__clkbuf_4 T22Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6286));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R0_INV_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6322));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R1_INV_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R2_INV_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R2_INV_1 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6358));
  sky130_fd_sc_hd__clkbuf_4 T22Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6394));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R0_INV_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6430));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R1_INV_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R2_INV_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R2_INV_1 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6466));
  sky130_fd_sc_hd__clkbuf_4 T22Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B563));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R0_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B599));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R1_INV_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R2_INV_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R2_INV_1 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B635));
  sky130_fd_sc_hd__clkbuf_4 T22Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6502));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R0_INV_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6538));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R1_INV_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R2_INV_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R2_INV_1 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6574));
  sky130_fd_sc_hd__clkbuf_4 T22Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6610));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R0_INV_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6646));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R1_INV_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R2_INV_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R2_INV_1 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6682));
  sky130_fd_sc_hd__clkbuf_4 T22Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6718));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R0_INV_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6754));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R1_INV_0 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R2_INV_0 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R2_INV_1 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6790));
  sky130_fd_sc_hd__clkbuf_4 T22Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6826));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R0_INV_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6862));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R1_INV_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R2_INV_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R2_INV_1 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6898));
  sky130_fd_sc_hd__clkbuf_4 T22Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6934));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R0_INV_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6970));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R1_INV_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R2_INV_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R2_INV_1 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7006));
  sky130_fd_sc_hd__clkbuf_4 T22Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7042));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R0_INV_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7078));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R1_INV_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R2_INV_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R2_INV_1 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7114));
  sky130_fd_sc_hd__clkbuf_4 T22Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7150));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R0_INV_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7186));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R1_INV_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R2_INV_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R2_INV_1 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7222));
  sky130_fd_sc_hd__clkbuf_4 T22Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7258));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R0_INV_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7294));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R1_INV_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R2_INV_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R2_INV_1 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7330));
  sky130_fd_sc_hd__clkbuf_4 T22Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7366));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R0_INV_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7402));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R1_INV_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R2_INV_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R2_INV_1 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7438));
  sky130_fd_sc_hd__clkbuf_4 T22Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7474));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R0_INV_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7510));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R1_INV_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R2_INV_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R2_INV_1 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7546));
  sky130_fd_sc_hd__clkbuf_4 T22Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B671));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R0_INV_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B707));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R1_INV_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R2_INV_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R2_INV_1 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B743));
  sky130_fd_sc_hd__clkbuf_4 T22Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7582));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R0_INV_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7618));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R1_INV_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R2_INV_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R2_INV_1 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7654));
  sky130_fd_sc_hd__clkbuf_4 T22Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7690));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R0_INV_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7726));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R1_INV_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R2_INV_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R2_INV_1 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7762));
  sky130_fd_sc_hd__clkbuf_4 T22Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7798));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R0_INV_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7834));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R1_INV_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R2_INV_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R2_INV_1 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7870));
  sky130_fd_sc_hd__clkbuf_4 T22Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7906));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R0_INV_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7942));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R1_INV_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R2_INV_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R2_INV_1 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7978));
  sky130_fd_sc_hd__clkbuf_4 T22Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8014));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R0_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8050));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R1_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R2_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R2_INV_1 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8086));
  sky130_fd_sc_hd__clkbuf_4 T22Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8122));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R0_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8158));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R1_INV_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R2_INV_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R2_INV_1 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8194));
  sky130_fd_sc_hd__clkbuf_4 T22Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8230));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R0_INV_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8266));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R1_INV_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R2_INV_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R2_INV_1 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8302));
  sky130_fd_sc_hd__clkbuf_4 T22Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8338));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R0_INV_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8374));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R1_INV_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R2_INV_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R2_INV_1 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8410));
  sky130_fd_sc_hd__clkbuf_4 T22Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8446));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R0_INV_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8482));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R1_INV_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R2_INV_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R2_INV_1 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8518));
  sky130_fd_sc_hd__clkbuf_4 T22Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8554));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R0_INV_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8590));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R1_INV_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R2_INV_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R2_INV_1 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8626));
  sky130_fd_sc_hd__clkbuf_4 T22Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B779));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R0_INV_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B815));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R1_INV_0 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R2_INV_0 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R2_INV_1 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B851));
  sky130_fd_sc_hd__clkbuf_4 T22Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8662));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R0_INV_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8698));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R1_INV_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R2_INV_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R2_INV_1 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8734));
  sky130_fd_sc_hd__clkbuf_4 T22Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8770));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R0_INV_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8806));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R1_INV_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R2_INV_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R2_INV_1 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8842));
  sky130_fd_sc_hd__clkbuf_4 T22Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8878));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R0_INV_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8914));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R1_INV_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R2_INV_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R2_INV_1 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8950));
  sky130_fd_sc_hd__clkbuf_4 T22Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8986));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R0_INV_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9022));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R1_INV_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R2_INV_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R2_INV_1 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9058));
  sky130_fd_sc_hd__clkbuf_4 T22Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9094));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R0_INV_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9130));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R1_INV_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R2_INV_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R2_INV_1 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9166));
  sky130_fd_sc_hd__clkbuf_4 T22Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9202));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R0_INV_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9238));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R1_INV_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R2_INV_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R2_INV_1 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9274));
  sky130_fd_sc_hd__clkbuf_4 T22Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9310));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R0_INV_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9346));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R1_INV_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R2_INV_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R2_INV_1 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9382));
  sky130_fd_sc_hd__clkbuf_4 T22Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9418));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R0_INV_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9454));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R1_INV_0 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R2_INV_0 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R2_INV_1 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9490));
  sky130_fd_sc_hd__clkbuf_4 T22Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9526));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R0_INV_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9562));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R1_INV_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R2_INV_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R2_INV_1 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9598));
  sky130_fd_sc_hd__clkbuf_4 T22Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9634));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R0_INV_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9670));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R1_INV_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R2_INV_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R2_INV_1 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9706));
  sky130_fd_sc_hd__clkbuf_4 T22Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B887));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R0_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B923));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R1_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R2_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R2_INV_1 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B959));
  sky130_fd_sc_hd__clkbuf_4 T22Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B995));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R0_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1031));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R1_INV_0 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R2_INV_0 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R2_INV_1 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1067));
  sky130_fd_sc_hd__clkbuf_4 T23Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B33));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R0_INV_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B68));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R1_INV_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R2_INV_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R2_INV_1 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B103));
  sky130_fd_sc_hd__clkbuf_4 T23Y10__R0_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B69));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R0_INV_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1140));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R1_INV_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R2_INV_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R2_INV_1 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1176));
  sky130_fd_sc_hd__clkbuf_4 T23Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1212));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R0_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y11__R1_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B78));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R1_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R2_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R2_INV_1 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1284));
  sky130_fd_sc_hd__clkbuf_4 T23Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1320));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R0_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1356));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R1_INV_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R2_INV_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R2_INV_1 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y12__R3_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B87));
  sky130_fd_sc_hd__clkbuf_4 T23Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1428));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R0_INV_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1464));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R1_INV_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R2_INV_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R2_INV_1 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1500));
  sky130_fd_sc_hd__clkbuf_4 T23Y14__R0_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B6));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R0_INV_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1571));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R1_INV_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R2_INV_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R2_INV_1 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1607));
  sky130_fd_sc_hd__clkbuf_4 T23Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1643));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R0_INV_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1679));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R1_INV_0 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R2_INV_0 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R2_INV_1 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1715));
  sky130_fd_sc_hd__clkbuf_4 T23Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1751));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R0_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1787));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R1_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R2_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R2_INV_1 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1823));
  sky130_fd_sc_hd__clkbuf_4 T23Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1859));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R0_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1895));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R1_INV_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R2_INV_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R2_INV_1 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1931));
  sky130_fd_sc_hd__clkbuf_4 T23Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1967));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R0_INV_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2003));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R1_INV_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R2_INV_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R2_INV_1 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2039));
  sky130_fd_sc_hd__clkbuf_4 T23Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2075));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R0_INV_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2111));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R1_INV_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R2_INV_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R2_INV_1 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2147));
  sky130_fd_sc_hd__clkbuf_4 T23Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B138));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R0_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B173));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R1_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R2_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R2_INV_1 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y1__R3_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B13));
  sky130_fd_sc_hd__clkbuf_4 T23Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2183));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R0_INV_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2219));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R1_INV_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R2_INV_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R2_INV_1 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2255));
  sky130_fd_sc_hd__clkbuf_4 T23Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2291));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R0_INV_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2327));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R1_INV_0 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R2_INV_0 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R2_INV_1 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2363));
  sky130_fd_sc_hd__clkbuf_4 T23Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2399));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R0_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2435));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R1_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R2_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R2_INV_1 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2471));
  sky130_fd_sc_hd__clkbuf_4 T23Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2507));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R0_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2543));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R1_INV_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R2_INV_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R2_INV_1 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2579));
  sky130_fd_sc_hd__clkbuf_4 T23Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2615));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R0_INV_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2651));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R1_INV_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R2_INV_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R2_INV_1 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2687));
  sky130_fd_sc_hd__clkbuf_4 T23Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2723));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R0_INV_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2759));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R1_INV_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R2_INV_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R2_INV_1 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2795));
  sky130_fd_sc_hd__clkbuf_4 T23Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2831));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R0_INV_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2867));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R1_INV_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R2_INV_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R2_INV_1 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2903));
  sky130_fd_sc_hd__clkbuf_4 T23Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2939));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R0_INV_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2975));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R1_INV_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R2_INV_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R2_INV_1 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3011));
  sky130_fd_sc_hd__clkbuf_4 T23Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3047));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R0_INV_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3083));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R1_INV_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R2_INV_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R2_INV_1 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3119));
  sky130_fd_sc_hd__clkbuf_4 T23Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3155));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R0_INV_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3191));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R1_INV_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R2_INV_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R2_INV_1 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3227));
  sky130_fd_sc_hd__clkbuf_4 T23Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B243));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R0_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B278));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R1_INV_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R2_INV_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R2_INV_1 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B314));
  sky130_fd_sc_hd__clkbuf_4 T23Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3263));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R0_INV_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3299));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R1_INV_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R2_INV_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R2_INV_1 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3335));
  sky130_fd_sc_hd__clkbuf_4 T23Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3371));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R0_INV_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3407));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R1_INV_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R2_INV_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R2_INV_1 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3443));
  sky130_fd_sc_hd__clkbuf_4 T23Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3479));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R0_INV_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3515));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R1_INV_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R2_INV_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R2_INV_1 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3551));
  sky130_fd_sc_hd__clkbuf_4 T23Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3587));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R0_INV_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3623));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R1_INV_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R2_INV_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R2_INV_1 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3659));
  sky130_fd_sc_hd__clkbuf_4 T23Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3695));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R0_INV_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3731));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R1_INV_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R2_INV_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R2_INV_1 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3767));
  sky130_fd_sc_hd__clkbuf_4 T23Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3803));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R0_INV_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3839));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R1_INV_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R2_INV_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R2_INV_1 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3875));
  sky130_fd_sc_hd__clkbuf_4 T23Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3911));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R0_INV_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3947));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R1_INV_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R2_INV_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R2_INV_1 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3983));
  sky130_fd_sc_hd__clkbuf_4 T23Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4019));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R0_INV_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4055));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R1_INV_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R2_INV_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R2_INV_1 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4091));
  sky130_fd_sc_hd__clkbuf_4 T23Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4127));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R0_INV_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4163));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R1_INV_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R2_INV_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R2_INV_1 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4199));
  sky130_fd_sc_hd__clkbuf_4 T23Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4235));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R0_INV_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4271));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R1_INV_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R2_INV_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R2_INV_1 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4307));
  sky130_fd_sc_hd__clkbuf_4 T23Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B349));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R0_INV_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y3__R1_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B24));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R1_INV_0 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R2_INV_0 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R2_INV_1 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B420));
  sky130_fd_sc_hd__clkbuf_4 T23Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4343));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R0_INV_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4379));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R1_INV_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R2_INV_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R2_INV_1 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4415));
  sky130_fd_sc_hd__clkbuf_4 T23Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4451));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R0_INV_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4487));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R1_INV_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R2_INV_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R2_INV_1 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4523));
  sky130_fd_sc_hd__clkbuf_4 T23Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4559));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R0_INV_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4595));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R1_INV_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R2_INV_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R2_INV_1 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4631));
  sky130_fd_sc_hd__clkbuf_4 T23Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4667));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R0_INV_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4703));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R1_INV_0 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R2_INV_0 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R2_INV_1 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4739));
  sky130_fd_sc_hd__clkbuf_4 T23Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4775));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R0_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4811));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R1_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R2_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R2_INV_1 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4847));
  sky130_fd_sc_hd__clkbuf_4 T23Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4883));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R0_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4919));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R1_INV_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R2_INV_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R2_INV_1 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4955));
  sky130_fd_sc_hd__clkbuf_4 T23Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4991));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R0_INV_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5027));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R1_INV_0 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R2_INV_0 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R2_INV_1 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5063));
  sky130_fd_sc_hd__clkbuf_4 T23Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5099));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R0_INV_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5135));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R1_INV_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R2_INV_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R2_INV_1 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5171));
  sky130_fd_sc_hd__clkbuf_4 T23Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5207));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R0_INV_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5243));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R1_INV_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R2_INV_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R2_INV_1 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5279));
  sky130_fd_sc_hd__clkbuf_4 T23Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5315));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R0_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5351));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R1_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R2_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R2_INV_1 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5387));
  sky130_fd_sc_hd__clkbuf_4 T23Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B456));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R0_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B492));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R1_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R2_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R2_INV_1 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y4__R3_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B33));
  sky130_fd_sc_hd__clkbuf_4 T23Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5423));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R0_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5459));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R1_INV_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R2_INV_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R2_INV_1 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5495));
  sky130_fd_sc_hd__clkbuf_4 T23Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5531));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R0_INV_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5567));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R1_INV_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R2_INV_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R2_INV_1 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5603));
  sky130_fd_sc_hd__clkbuf_4 T23Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5639));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R0_INV_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5675));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R1_INV_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R2_INV_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R2_INV_1 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5711));
  sky130_fd_sc_hd__clkbuf_4 T23Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5747));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R0_INV_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5783));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R1_INV_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R2_INV_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R2_INV_1 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5819));
  sky130_fd_sc_hd__clkbuf_4 T23Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5855));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R0_INV_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5891));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R1_INV_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R2_INV_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R2_INV_1 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5927));
  sky130_fd_sc_hd__clkbuf_4 T23Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5963));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R0_INV_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5999));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R1_INV_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R2_INV_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R2_INV_1 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6035));
  sky130_fd_sc_hd__clkbuf_4 T23Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6071));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R0_INV_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6107));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R1_INV_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R2_INV_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R2_INV_1 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6143));
  sky130_fd_sc_hd__clkbuf_4 T23Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6179));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R0_INV_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6215));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R1_INV_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R2_INV_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R2_INV_1 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6251));
  sky130_fd_sc_hd__clkbuf_4 T23Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6287));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R0_INV_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6323));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R1_INV_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R2_INV_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R2_INV_1 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6359));
  sky130_fd_sc_hd__clkbuf_4 T23Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6395));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R0_INV_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6431));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R1_INV_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R2_INV_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R2_INV_1 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6467));
  sky130_fd_sc_hd__clkbuf_4 T23Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B564));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R0_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B600));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R1_INV_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R2_INV_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R2_INV_1 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B636));
  sky130_fd_sc_hd__clkbuf_4 T23Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6503));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R0_INV_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6539));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R1_INV_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R2_INV_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R2_INV_1 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6575));
  sky130_fd_sc_hd__clkbuf_4 T23Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6611));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R0_INV_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6647));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R1_INV_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R2_INV_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R2_INV_1 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6683));
  sky130_fd_sc_hd__clkbuf_4 T23Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6719));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R0_INV_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6755));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R1_INV_0 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R2_INV_0 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R2_INV_1 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6791));
  sky130_fd_sc_hd__clkbuf_4 T23Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6827));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R0_INV_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6863));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R1_INV_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R2_INV_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R2_INV_1 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6899));
  sky130_fd_sc_hd__clkbuf_4 T23Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6935));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R0_INV_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6971));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R1_INV_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R2_INV_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R2_INV_1 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B7007));
  sky130_fd_sc_hd__clkbuf_4 T23Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7043));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R0_INV_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7079));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R1_INV_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R2_INV_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R2_INV_1 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7115));
  sky130_fd_sc_hd__clkbuf_4 T23Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7151));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R0_INV_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7187));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R1_INV_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R2_INV_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R2_INV_1 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7223));
  sky130_fd_sc_hd__clkbuf_4 T23Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7259));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R0_INV_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7295));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R1_INV_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R2_INV_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R2_INV_1 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7331));
  sky130_fd_sc_hd__clkbuf_4 T23Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7367));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R0_INV_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7403));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R1_INV_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R2_INV_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R2_INV_1 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7439));
  sky130_fd_sc_hd__clkbuf_4 T23Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7475));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R0_INV_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7511));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R1_INV_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R2_INV_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R2_INV_1 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7547));
  sky130_fd_sc_hd__clkbuf_4 T23Y6__R0_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B42));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R0_INV_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B708));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R1_INV_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R2_INV_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R2_INV_1 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B744));
  sky130_fd_sc_hd__clkbuf_4 T23Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7583));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R0_INV_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7619));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R1_INV_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R2_INV_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R2_INV_1 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7655));
  sky130_fd_sc_hd__clkbuf_4 T23Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7691));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R0_INV_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7727));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R1_INV_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R2_INV_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R2_INV_1 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7763));
  sky130_fd_sc_hd__clkbuf_4 T23Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7799));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R0_INV_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7835));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R1_INV_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R2_INV_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R2_INV_1 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7871));
  sky130_fd_sc_hd__clkbuf_4 T23Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7907));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R0_INV_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7943));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R1_INV_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R2_INV_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R2_INV_1 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7979));
  sky130_fd_sc_hd__clkbuf_4 T23Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8015));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R0_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8051));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R1_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R2_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R2_INV_1 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8087));
  sky130_fd_sc_hd__clkbuf_4 T23Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8123));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R0_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8159));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R1_INV_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R2_INV_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R2_INV_1 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8195));
  sky130_fd_sc_hd__clkbuf_4 T23Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8231));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R0_INV_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8267));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R1_INV_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R2_INV_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R2_INV_1 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8303));
  sky130_fd_sc_hd__clkbuf_4 T23Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8339));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R0_INV_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8375));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R1_INV_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R2_INV_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R2_INV_1 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8411));
  sky130_fd_sc_hd__clkbuf_4 T23Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8447));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R0_INV_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8483));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R1_INV_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R2_INV_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R2_INV_1 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8519));
  sky130_fd_sc_hd__clkbuf_4 T23Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8555));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R0_INV_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8591));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R1_INV_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R2_INV_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R2_INV_1 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8627));
  sky130_fd_sc_hd__clkbuf_4 T23Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B780));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R0_INV_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y7__R1_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B51));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R1_INV_0 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R2_INV_0 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R2_INV_1 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B852));
  sky130_fd_sc_hd__clkbuf_4 T23Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8663));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R0_INV_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8699));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R1_INV_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R2_INV_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R2_INV_1 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8735));
  sky130_fd_sc_hd__clkbuf_4 T23Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8771));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R0_INV_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8807));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R1_INV_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R2_INV_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R2_INV_1 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8843));
  sky130_fd_sc_hd__clkbuf_4 T23Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8879));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R0_INV_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8915));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R1_INV_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R2_INV_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R2_INV_1 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8951));
  sky130_fd_sc_hd__clkbuf_4 T23Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8987));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R0_INV_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9023));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R1_INV_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R2_INV_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R2_INV_1 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9059));
  sky130_fd_sc_hd__clkbuf_4 T23Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9095));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R0_INV_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9131));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R1_INV_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R2_INV_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R2_INV_1 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9167));
  sky130_fd_sc_hd__clkbuf_4 T23Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9203));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R0_INV_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9239));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R1_INV_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R2_INV_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R2_INV_1 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9275));
  sky130_fd_sc_hd__clkbuf_4 T23Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9311));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R0_INV_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9347));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R1_INV_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R2_INV_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R2_INV_1 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9383));
  sky130_fd_sc_hd__clkbuf_4 T23Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9419));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R0_INV_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9455));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R1_INV_0 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R2_INV_0 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R2_INV_1 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9491));
  sky130_fd_sc_hd__clkbuf_4 T23Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9527));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R0_INV_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9563));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R1_INV_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R2_INV_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R2_INV_1 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9599));
  sky130_fd_sc_hd__clkbuf_4 T23Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9635));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R0_INV_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9671));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R1_INV_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R2_INV_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R2_INV_1 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9707));
  sky130_fd_sc_hd__clkbuf_4 T23Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B888));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R0_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B924));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R1_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R2_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R2_INV_1 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y8__R3_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B60));
  sky130_fd_sc_hd__clkbuf_4 T23Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B996));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R0_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1032));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R1_INV_0 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R2_INV_0 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R2_INV_1 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1068));
  sky130_fd_sc_hd__clkbuf_4 T24Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B34));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R0_INV_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B69));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R1_INV_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R2_INV_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R2_INV_1 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B104));
  sky130_fd_sc_hd__clkbuf_4 T24Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1105));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R0_INV_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1141));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R1_INV_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R2_INV_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R2_INV_1 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1177));
  sky130_fd_sc_hd__clkbuf_4 T24Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1213));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R0_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1249));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R1_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R2_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R2_INV_1 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1285));
  sky130_fd_sc_hd__clkbuf_4 T24Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1321));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R0_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1357));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R1_INV_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R2_INV_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R2_INV_1 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1393));
  sky130_fd_sc_hd__clkbuf_4 T24Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1429));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R0_INV_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1465));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R1_INV_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R2_INV_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R2_INV_1 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1501));
  sky130_fd_sc_hd__clkbuf_4 T24Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1537));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R0_INV_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1572));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R1_INV_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R2_INV_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R2_INV_1 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1608));
  sky130_fd_sc_hd__clkbuf_4 T24Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1644));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R0_INV_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y15__R1_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B105));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R1_INV_0 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R2_INV_0 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R2_INV_1 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1716));
  sky130_fd_sc_hd__clkbuf_4 T24Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1752));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R0_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1788));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R1_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R2_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R2_INV_1 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y16__R3_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B114));
  sky130_fd_sc_hd__clkbuf_4 T24Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1860));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R0_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1896));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R1_INV_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R2_INV_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R2_INV_1 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1932));
  sky130_fd_sc_hd__clkbuf_4 T24Y18__R0_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B123));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R0_INV_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2004));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R1_INV_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R2_INV_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R2_INV_1 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2040));
  sky130_fd_sc_hd__clkbuf_4 T24Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2076));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R0_INV_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y19__R1_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B132));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R1_INV_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R2_INV_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R2_INV_1 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2148));
  sky130_fd_sc_hd__clkbuf_4 T24Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B139));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R0_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B174));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R1_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R2_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R2_INV_1 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B209));
  sky130_fd_sc_hd__clkbuf_4 T24Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2184));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R0_INV_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2220));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R1_INV_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R2_INV_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R2_INV_1 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y20__R3_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B141));
  sky130_fd_sc_hd__clkbuf_4 T24Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2292));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R0_INV_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2328));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R1_INV_0 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R2_INV_0 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R2_INV_1 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2364));
  sky130_fd_sc_hd__clkbuf_4 T24Y22__R0_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B150));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R0_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2436));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R1_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R2_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R2_INV_1 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2472));
  sky130_fd_sc_hd__clkbuf_4 T24Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2508));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R0_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y23__R1_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B159));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R1_INV_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R2_INV_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R2_INV_1 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2580));
  sky130_fd_sc_hd__clkbuf_4 T24Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2616));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R0_INV_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2652));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R1_INV_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R2_INV_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R2_INV_1 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y24__R3_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B168));
  sky130_fd_sc_hd__clkbuf_4 T24Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2724));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R0_INV_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2760));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R1_INV_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R2_INV_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R2_INV_1 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2796));
  sky130_fd_sc_hd__clkbuf_4 T24Y26__R0_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B177));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R0_INV_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2868));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R1_INV_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R2_INV_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R2_INV_1 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2904));
  sky130_fd_sc_hd__clkbuf_4 T24Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2940));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R0_INV_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y27__R1_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B186));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R1_INV_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R2_INV_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R2_INV_1 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3012));
  sky130_fd_sc_hd__clkbuf_4 T24Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3048));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R0_INV_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3084));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R1_INV_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R2_INV_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R2_INV_1 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y28__R3_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B195));
  sky130_fd_sc_hd__clkbuf_4 T24Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3156));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R0_INV_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3192));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R1_INV_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R2_INV_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R2_INV_1 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3228));
  sky130_fd_sc_hd__clkbuf_4 T24Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B244));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R0_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B279));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R1_INV_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R2_INV_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R2_INV_1 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B315));
  sky130_fd_sc_hd__clkbuf_4 T24Y30__R0_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B204));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R0_INV_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3300));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R1_INV_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R2_INV_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R2_INV_1 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3336));
  sky130_fd_sc_hd__clkbuf_4 T24Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3372));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R0_INV_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y31__R1_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B213));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R1_INV_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R2_INV_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R2_INV_1 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3444));
  sky130_fd_sc_hd__clkbuf_4 T24Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3480));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R0_INV_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3516));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R1_INV_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R2_INV_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R2_INV_1 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y32__R3_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B222));
  sky130_fd_sc_hd__clkbuf_4 T24Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3588));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R0_INV_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3624));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R1_INV_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R2_INV_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R2_INV_1 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3660));
  sky130_fd_sc_hd__clkbuf_4 T24Y34__R0_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B231));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R0_INV_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3732));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R1_INV_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R2_INV_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R2_INV_1 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3768));
  sky130_fd_sc_hd__clkbuf_4 T24Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3804));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R0_INV_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y35__R1_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B15));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R1_INV_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R2_INV_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R2_INV_1 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3876));
  sky130_fd_sc_hd__clkbuf_4 T24Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3912));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R0_INV_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3948));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R1_INV_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R2_INV_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R2_INV_1 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y36__R3_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B249));
  sky130_fd_sc_hd__clkbuf_4 T24Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4020));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R0_INV_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4056));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R1_INV_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R2_INV_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R2_INV_1 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4092));
  sky130_fd_sc_hd__clkbuf_4 T24Y38__R0_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B258));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R0_INV_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4164));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R1_INV_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R2_INV_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R2_INV_1 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4200));
  sky130_fd_sc_hd__clkbuf_4 T24Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4236));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R0_INV_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y39__R1_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B267));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R1_INV_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R2_INV_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R2_INV_1 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4308));
  sky130_fd_sc_hd__clkbuf_4 T24Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B350));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R0_INV_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B385));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R1_INV_0 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R2_INV_0 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R2_INV_1 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B421));
  sky130_fd_sc_hd__clkbuf_4 T24Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4344));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R0_INV_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4380));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R1_INV_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R2_INV_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R2_INV_1 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y40__R3_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B276));
  sky130_fd_sc_hd__clkbuf_4 T24Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4452));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R0_INV_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4488));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R1_INV_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R2_INV_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R2_INV_1 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4524));
  sky130_fd_sc_hd__clkbuf_4 T24Y42__R0_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B285));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R0_INV_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4596));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R1_INV_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R2_INV_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R2_INV_1 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4632));
  sky130_fd_sc_hd__clkbuf_4 T24Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4668));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R0_INV_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y43__R1_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B294));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R1_INV_0 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R2_INV_0 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R2_INV_1 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4740));
  sky130_fd_sc_hd__clkbuf_4 T24Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4776));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R0_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4812));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R1_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R2_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R2_INV_1 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y44__R3_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B303));
  sky130_fd_sc_hd__clkbuf_4 T24Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4884));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R0_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4920));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R1_INV_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R2_INV_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R2_INV_1 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4956));
  sky130_fd_sc_hd__clkbuf_4 T24Y46__R0_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B312));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R0_INV_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5028));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R1_INV_0 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R2_INV_0 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R2_INV_1 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5064));
  sky130_fd_sc_hd__clkbuf_4 T24Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5100));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R0_INV_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y47__R1_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B321));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R1_INV_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R2_INV_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R2_INV_1 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5172));
  sky130_fd_sc_hd__clkbuf_4 T24Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5208));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R0_INV_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5244));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R1_INV_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R2_INV_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R2_INV_1 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y48__R3_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B330));
  sky130_fd_sc_hd__clkbuf_4 T24Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5316));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R0_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5352));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R1_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R2_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R2_INV_1 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5388));
  sky130_fd_sc_hd__clkbuf_4 T24Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B457));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R0_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B493));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R1_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R2_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R2_INV_1 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B529));
  sky130_fd_sc_hd__clkbuf_4 T24Y50__R0_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B339));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R0_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5460));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R1_INV_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R2_INV_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R2_INV_1 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5496));
  sky130_fd_sc_hd__clkbuf_4 T24Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5532));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R0_INV_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y51__R1_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B348));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R1_INV_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R2_INV_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R2_INV_1 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5604));
  sky130_fd_sc_hd__clkbuf_4 T24Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5640));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R0_INV_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5676));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R1_INV_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R2_INV_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R2_INV_1 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y52__R3_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B357));
  sky130_fd_sc_hd__clkbuf_4 T24Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5748));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R0_INV_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5784));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R1_INV_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R2_INV_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R2_INV_1 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5820));
  sky130_fd_sc_hd__clkbuf_4 T24Y54__R0_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B366));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R0_INV_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5892));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R1_INV_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R2_INV_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R2_INV_1 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5928));
  sky130_fd_sc_hd__clkbuf_4 T24Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5964));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R0_INV_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y55__R1_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B375));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R1_INV_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R2_INV_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R2_INV_1 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6036));
  sky130_fd_sc_hd__clkbuf_4 T24Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6072));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R0_INV_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6108));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R1_INV_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R2_INV_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R2_INV_1 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y56__R3_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B24));
  sky130_fd_sc_hd__clkbuf_4 T24Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6180));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R0_INV_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6216));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R1_INV_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R2_INV_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R2_INV_1 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6252));
  sky130_fd_sc_hd__clkbuf_4 T24Y58__R0_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B393));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R0_INV_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6324));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R1_INV_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R2_INV_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R2_INV_1 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6360));
  sky130_fd_sc_hd__clkbuf_4 T24Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6396));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R0_INV_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y59__R1_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B402));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R1_INV_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R2_INV_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R2_INV_1 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6468));
  sky130_fd_sc_hd__clkbuf_4 T24Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B565));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R0_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B601));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R1_INV_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R2_INV_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R2_INV_1 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B637));
  sky130_fd_sc_hd__clkbuf_4 T24Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6504));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R0_INV_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6540));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R1_INV_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R2_INV_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R2_INV_1 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y60__R3_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B411));
  sky130_fd_sc_hd__clkbuf_4 T24Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6612));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R0_INV_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6648));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R1_INV_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R2_INV_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R2_INV_1 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6684));
  sky130_fd_sc_hd__clkbuf_4 T24Y62__R0_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B420));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R0_INV_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6756));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R1_INV_0 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R2_INV_0 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R2_INV_1 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6792));
  sky130_fd_sc_hd__clkbuf_4 T24Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6828));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R0_INV_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y63__R1_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B429));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R1_INV_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R2_INV_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R2_INV_1 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6900));
  sky130_fd_sc_hd__clkbuf_4 T24Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6936));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R0_INV_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6972));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R1_INV_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R2_INV_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R2_INV_1 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y64__R3_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B438));
  sky130_fd_sc_hd__clkbuf_4 T24Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7044));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R0_INV_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7080));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R1_INV_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R2_INV_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R2_INV_1 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7116));
  sky130_fd_sc_hd__clkbuf_4 T24Y66__R0_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B447));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R0_INV_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7188));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R1_INV_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R2_INV_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R2_INV_1 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7224));
  sky130_fd_sc_hd__clkbuf_4 T24Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7260));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R0_INV_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y67__R1_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B456));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R1_INV_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R2_INV_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R2_INV_1 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7332));
  sky130_fd_sc_hd__clkbuf_4 T24Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7368));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R0_INV_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7404));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R1_INV_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R2_INV_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R2_INV_1 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y68__R3_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B465));
  sky130_fd_sc_hd__clkbuf_4 T24Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7476));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R0_INV_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7512));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R1_INV_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R2_INV_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R2_INV_1 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7548));
  sky130_fd_sc_hd__clkbuf_4 T24Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B673));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R0_INV_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B709));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R1_INV_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R2_INV_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R2_INV_1 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B745));
  sky130_fd_sc_hd__clkbuf_4 T24Y70__R0_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B474));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R0_INV_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7620));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R1_INV_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R2_INV_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R2_INV_1 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7656));
  sky130_fd_sc_hd__clkbuf_4 T24Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7692));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R0_INV_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y71__R1_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B483));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R1_INV_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R2_INV_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R2_INV_1 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7764));
  sky130_fd_sc_hd__clkbuf_4 T24Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7800));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R0_INV_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7836));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R1_INV_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R2_INV_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R2_INV_1 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y72__R3_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B492));
  sky130_fd_sc_hd__clkbuf_4 T24Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7908));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R0_INV_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7944));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R1_INV_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R2_INV_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R2_INV_1 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7980));
  sky130_fd_sc_hd__clkbuf_4 T24Y74__R0_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B501));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R0_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8052));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R1_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R2_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R2_INV_1 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8088));
  sky130_fd_sc_hd__clkbuf_4 T24Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8124));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R0_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y75__R1_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B510));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R1_INV_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R2_INV_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R2_INV_1 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8196));
  sky130_fd_sc_hd__clkbuf_4 T24Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8232));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R0_INV_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8268));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R1_INV_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R2_INV_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R2_INV_1 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y76__R3_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B519));
  sky130_fd_sc_hd__clkbuf_4 T24Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8340));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R0_INV_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8376));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R1_INV_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R2_INV_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R2_INV_1 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8412));
  sky130_fd_sc_hd__clkbuf_4 T24Y78__R0_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B33));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R0_INV_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8484));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R1_INV_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R2_INV_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R2_INV_1 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8520));
  sky130_fd_sc_hd__clkbuf_4 T24Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8556));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R0_INV_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y79__R1_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B537));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R1_INV_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R2_INV_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R2_INV_1 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8628));
  sky130_fd_sc_hd__clkbuf_4 T24Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B781));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R0_INV_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B817));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R1_INV_0 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R2_INV_0 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R2_INV_1 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B853));
  sky130_fd_sc_hd__clkbuf_4 T24Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8664));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R0_INV_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8700));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R1_INV_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R2_INV_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R2_INV_1 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y80__R3_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B546));
  sky130_fd_sc_hd__clkbuf_4 T24Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8772));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R0_INV_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8808));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R1_INV_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R2_INV_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R2_INV_1 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8844));
  sky130_fd_sc_hd__clkbuf_4 T24Y82__R0_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B555));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R0_INV_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8916));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R1_INV_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R2_INV_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R2_INV_1 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8952));
  sky130_fd_sc_hd__clkbuf_4 T24Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8988));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R0_INV_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y83__R1_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B564));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R1_INV_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R2_INV_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R2_INV_1 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9060));
  sky130_fd_sc_hd__clkbuf_4 T24Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9096));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R0_INV_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9132));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R1_INV_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R2_INV_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R2_INV_1 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y84__R3_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B573));
  sky130_fd_sc_hd__clkbuf_4 T24Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9204));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R0_INV_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9240));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R1_INV_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R2_INV_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R2_INV_1 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9276));
  sky130_fd_sc_hd__clkbuf_4 T24Y86__R0_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B582));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R0_INV_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9348));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R1_INV_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R2_INV_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R2_INV_1 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9384));
  sky130_fd_sc_hd__clkbuf_4 T24Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9420));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R0_INV_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y87__R1_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B591));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R1_INV_0 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R2_INV_0 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R2_INV_1 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9492));
  sky130_fd_sc_hd__clkbuf_4 T24Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9528));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R0_INV_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9564));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R1_INV_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R2_INV_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R2_INV_1 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y88__R3_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B600));
  sky130_fd_sc_hd__clkbuf_4 T24Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9636));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R0_INV_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9672));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R1_INV_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R2_INV_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R2_INV_1 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9708));
  sky130_fd_sc_hd__clkbuf_4 T24Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B889));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R0_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B925));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R1_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R2_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R2_INV_1 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B961));
  sky130_fd_sc_hd__clkbuf_4 T24Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B997));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R0_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1033));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R1_INV_0 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R2_INV_0 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R2_INV_1 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1069));
  sky130_fd_sc_hd__clkbuf_4 T25Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B35));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R0_INV_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B70));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R1_INV_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R2_INV_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R2_INV_1 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B105));
  sky130_fd_sc_hd__clkbuf_4 T25Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1106));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R0_INV_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1142));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R1_INV_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R2_INV_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R2_INV_1 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1178));
  sky130_fd_sc_hd__clkbuf_4 T25Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1214));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R0_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1250));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R1_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R2_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R2_INV_1 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1286));
  sky130_fd_sc_hd__clkbuf_4 T25Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1322));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R0_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1358));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R1_INV_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R2_INV_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R2_INV_1 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1394));
  sky130_fd_sc_hd__clkbuf_4 T25Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1430));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R0_INV_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1466));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R1_INV_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R2_INV_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R2_INV_1 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1502));
  sky130_fd_sc_hd__clkbuf_4 T25Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1538));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R0_INV_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1573));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R1_INV_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R2_INV_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R2_INV_1 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1609));
  sky130_fd_sc_hd__clkbuf_4 T25Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1645));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R0_INV_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1681));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R1_INV_0 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R2_INV_0 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R2_INV_1 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1717));
  sky130_fd_sc_hd__clkbuf_4 T25Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1753));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R0_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1789));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R1_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R2_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R2_INV_1 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1825));
  sky130_fd_sc_hd__clkbuf_4 T25Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1861));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R0_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1897));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R1_INV_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R2_INV_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R2_INV_1 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1933));
  sky130_fd_sc_hd__clkbuf_4 T25Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1969));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R0_INV_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2005));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R1_INV_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R2_INV_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R2_INV_1 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2041));
  sky130_fd_sc_hd__clkbuf_4 T25Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2077));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R0_INV_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2113));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R1_INV_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R2_INV_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R2_INV_1 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2149));
  sky130_fd_sc_hd__clkbuf_4 T25Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B140));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R0_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y1__R1_BUF_0 (.A(clk_L1_B10), .X(clk_L0_B175));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R1_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R2_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R2_INV_1 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B210));
  sky130_fd_sc_hd__clkbuf_4 T25Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2185));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R0_INV_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2221));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R1_INV_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R2_INV_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R2_INV_1 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2257));
  sky130_fd_sc_hd__clkbuf_4 T25Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2293));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R0_INV_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2329));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R1_INV_0 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R2_INV_0 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R2_INV_1 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2365));
  sky130_fd_sc_hd__clkbuf_4 T25Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2401));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R0_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2437));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R1_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R2_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R2_INV_1 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2473));
  sky130_fd_sc_hd__clkbuf_4 T25Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2509));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R0_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2545));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R1_INV_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R2_INV_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R2_INV_1 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2581));
  sky130_fd_sc_hd__clkbuf_4 T25Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2617));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R0_INV_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2653));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R1_INV_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R2_INV_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R2_INV_1 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2689));
  sky130_fd_sc_hd__clkbuf_4 T25Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2725));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R0_INV_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2761));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R1_INV_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R2_INV_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R2_INV_1 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2797));
  sky130_fd_sc_hd__clkbuf_4 T25Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2833));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R0_INV_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2869));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R1_INV_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R2_INV_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R2_INV_1 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2905));
  sky130_fd_sc_hd__clkbuf_4 T25Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2941));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R0_INV_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2977));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R1_INV_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R2_INV_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R2_INV_1 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3013));
  sky130_fd_sc_hd__clkbuf_4 T25Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3049));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R0_INV_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3085));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R1_INV_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R2_INV_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R2_INV_1 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3121));
  sky130_fd_sc_hd__clkbuf_4 T25Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3157));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R0_INV_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3193));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R1_INV_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R2_INV_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R2_INV_1 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3229));
  sky130_fd_sc_hd__clkbuf_4 T25Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B245));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R0_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B280));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R1_INV_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R2_INV_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R2_INV_1 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B316));
  sky130_fd_sc_hd__clkbuf_4 T25Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3265));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R0_INV_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3301));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R1_INV_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R2_INV_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R2_INV_1 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3337));
  sky130_fd_sc_hd__clkbuf_4 T25Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3373));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R0_INV_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3409));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R1_INV_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R2_INV_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R2_INV_1 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3445));
  sky130_fd_sc_hd__clkbuf_4 T25Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3481));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R0_INV_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3517));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R1_INV_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R2_INV_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R2_INV_1 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3553));
  sky130_fd_sc_hd__clkbuf_4 T25Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3589));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R0_INV_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3625));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R1_INV_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R2_INV_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R2_INV_1 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3661));
  sky130_fd_sc_hd__clkbuf_4 T25Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3697));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R0_INV_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3733));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R1_INV_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R2_INV_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R2_INV_1 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3769));
  sky130_fd_sc_hd__clkbuf_4 T25Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3805));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R0_INV_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3841));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R1_INV_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R2_INV_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R2_INV_1 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3877));
  sky130_fd_sc_hd__clkbuf_4 T25Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3913));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R0_INV_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3949));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R1_INV_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R2_INV_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R2_INV_1 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3985));
  sky130_fd_sc_hd__clkbuf_4 T25Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4021));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R0_INV_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4057));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R1_INV_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R2_INV_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R2_INV_1 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4093));
  sky130_fd_sc_hd__clkbuf_4 T25Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4129));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R0_INV_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4165));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R1_INV_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R2_INV_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R2_INV_1 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4201));
  sky130_fd_sc_hd__clkbuf_4 T25Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4237));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R0_INV_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4273));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R1_INV_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R2_INV_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R2_INV_1 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4309));
  sky130_fd_sc_hd__clkbuf_4 T25Y3__R0_BUF_0 (.A(clk_L1_B21), .X(clk_L0_B351));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R0_INV_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B386));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R1_INV_0 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R2_INV_0 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R2_INV_1 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B422));
  sky130_fd_sc_hd__clkbuf_4 T25Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4345));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R0_INV_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4381));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R1_INV_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R2_INV_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R2_INV_1 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4417));
  sky130_fd_sc_hd__clkbuf_4 T25Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4453));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R0_INV_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4489));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R1_INV_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R2_INV_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R2_INV_1 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4525));
  sky130_fd_sc_hd__clkbuf_4 T25Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4561));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R0_INV_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4597));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R1_INV_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R2_INV_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R2_INV_1 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4633));
  sky130_fd_sc_hd__clkbuf_4 T25Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4669));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R0_INV_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4705));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R1_INV_0 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R2_INV_0 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R2_INV_1 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4741));
  sky130_fd_sc_hd__clkbuf_4 T25Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4777));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R0_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4813));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R1_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R2_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R2_INV_1 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4849));
  sky130_fd_sc_hd__clkbuf_4 T25Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4885));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R0_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4921));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R1_INV_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R2_INV_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R2_INV_1 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4957));
  sky130_fd_sc_hd__clkbuf_4 T25Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4993));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R0_INV_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5029));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R1_INV_0 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R2_INV_0 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R2_INV_1 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5065));
  sky130_fd_sc_hd__clkbuf_4 T25Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5101));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R0_INV_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5137));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R1_INV_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R2_INV_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R2_INV_1 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5173));
  sky130_fd_sc_hd__clkbuf_4 T25Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5209));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R0_INV_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5245));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R1_INV_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R2_INV_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R2_INV_1 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5281));
  sky130_fd_sc_hd__clkbuf_4 T25Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5317));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R0_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5353));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R1_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R2_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R2_INV_1 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5389));
  sky130_fd_sc_hd__clkbuf_4 T25Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B458));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R0_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B494));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R1_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R2_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R2_INV_1 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B530));
  sky130_fd_sc_hd__clkbuf_4 T25Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5425));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R0_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5461));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R1_INV_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R2_INV_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R2_INV_1 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5497));
  sky130_fd_sc_hd__clkbuf_4 T25Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5533));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R0_INV_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5569));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R1_INV_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R2_INV_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R2_INV_1 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5605));
  sky130_fd_sc_hd__clkbuf_4 T25Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5641));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R0_INV_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5677));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R1_INV_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R2_INV_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R2_INV_1 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5713));
  sky130_fd_sc_hd__clkbuf_4 T25Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5749));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R0_INV_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5785));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R1_INV_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R2_INV_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R2_INV_1 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5821));
  sky130_fd_sc_hd__clkbuf_4 T25Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5857));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R0_INV_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5893));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R1_INV_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R2_INV_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R2_INV_1 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5929));
  sky130_fd_sc_hd__clkbuf_4 T25Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5965));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R0_INV_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6001));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R1_INV_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R2_INV_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R2_INV_1 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6037));
  sky130_fd_sc_hd__clkbuf_4 T25Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6073));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R0_INV_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6109));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R1_INV_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R2_INV_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R2_INV_1 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6145));
  sky130_fd_sc_hd__clkbuf_4 T25Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6181));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R0_INV_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6217));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R1_INV_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R2_INV_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R2_INV_1 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6253));
  sky130_fd_sc_hd__clkbuf_4 T25Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6289));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R0_INV_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6325));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R1_INV_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R2_INV_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R2_INV_1 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6361));
  sky130_fd_sc_hd__clkbuf_4 T25Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6397));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R0_INV_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6433));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R1_INV_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R2_INV_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R2_INV_1 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6469));
  sky130_fd_sc_hd__clkbuf_4 T25Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B566));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R0_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B602));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R1_INV_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R2_INV_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R2_INV_1 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B638));
  sky130_fd_sc_hd__clkbuf_4 T25Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6505));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R0_INV_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6541));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R1_INV_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R2_INV_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R2_INV_1 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6577));
  sky130_fd_sc_hd__clkbuf_4 T25Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6613));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R0_INV_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6649));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R1_INV_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R2_INV_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R2_INV_1 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6685));
  sky130_fd_sc_hd__clkbuf_4 T25Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6721));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R0_INV_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6757));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R1_INV_0 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R2_INV_0 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R2_INV_1 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6793));
  sky130_fd_sc_hd__clkbuf_4 T25Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6829));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R0_INV_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6865));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R1_INV_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R2_INV_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R2_INV_1 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6901));
  sky130_fd_sc_hd__clkbuf_4 T25Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6937));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R0_INV_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6973));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R1_INV_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R2_INV_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R2_INV_1 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7009));
  sky130_fd_sc_hd__clkbuf_4 T25Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7045));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R0_INV_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7081));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R1_INV_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R2_INV_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R2_INV_1 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7117));
  sky130_fd_sc_hd__clkbuf_4 T25Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7153));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R0_INV_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7189));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R1_INV_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R2_INV_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R2_INV_1 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7225));
  sky130_fd_sc_hd__clkbuf_4 T25Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7261));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R0_INV_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7297));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R1_INV_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R2_INV_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R2_INV_1 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7333));
  sky130_fd_sc_hd__clkbuf_4 T25Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7369));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R0_INV_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7405));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R1_INV_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R2_INV_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R2_INV_1 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7441));
  sky130_fd_sc_hd__clkbuf_4 T25Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7477));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R0_INV_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7513));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R1_INV_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R2_INV_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R2_INV_1 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7549));
  sky130_fd_sc_hd__clkbuf_4 T25Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B674));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R0_INV_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B710));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R1_INV_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R2_INV_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R2_INV_1 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B746));
  sky130_fd_sc_hd__clkbuf_4 T25Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7585));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R0_INV_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7621));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R1_INV_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R2_INV_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R2_INV_1 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7657));
  sky130_fd_sc_hd__clkbuf_4 T25Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7693));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R0_INV_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7729));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R1_INV_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R2_INV_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R2_INV_1 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7765));
  sky130_fd_sc_hd__clkbuf_4 T25Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7801));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R0_INV_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7837));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R1_INV_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R2_INV_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R2_INV_1 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7873));
  sky130_fd_sc_hd__clkbuf_4 T25Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7909));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R0_INV_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7945));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R1_INV_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R2_INV_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R2_INV_1 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7981));
  sky130_fd_sc_hd__clkbuf_4 T25Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8017));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R0_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8053));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R1_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R2_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R2_INV_1 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8089));
  sky130_fd_sc_hd__clkbuf_4 T25Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8125));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R0_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8161));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R1_INV_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R2_INV_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R2_INV_1 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8197));
  sky130_fd_sc_hd__clkbuf_4 T25Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8233));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R0_INV_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8269));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R1_INV_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R2_INV_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R2_INV_1 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8305));
  sky130_fd_sc_hd__clkbuf_4 T25Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8341));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R0_INV_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8377));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R1_INV_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R2_INV_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R2_INV_1 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8413));
  sky130_fd_sc_hd__clkbuf_4 T25Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8449));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R0_INV_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8485));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R1_INV_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R2_INV_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R2_INV_1 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8521));
  sky130_fd_sc_hd__clkbuf_4 T25Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8557));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R0_INV_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8593));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R1_INV_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R2_INV_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R2_INV_1 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8629));
  sky130_fd_sc_hd__clkbuf_4 T25Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B782));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R0_INV_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B818));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R1_INV_0 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R2_INV_0 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R2_INV_1 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B854));
  sky130_fd_sc_hd__clkbuf_4 T25Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8665));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R0_INV_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8701));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R1_INV_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R2_INV_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R2_INV_1 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8737));
  sky130_fd_sc_hd__clkbuf_4 T25Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8773));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R0_INV_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8809));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R1_INV_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R2_INV_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R2_INV_1 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8845));
  sky130_fd_sc_hd__clkbuf_4 T25Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8881));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R0_INV_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8917));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R1_INV_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R2_INV_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R2_INV_1 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8953));
  sky130_fd_sc_hd__clkbuf_4 T25Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8989));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R0_INV_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9025));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R1_INV_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R2_INV_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R2_INV_1 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9061));
  sky130_fd_sc_hd__clkbuf_4 T25Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9097));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R0_INV_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9133));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R1_INV_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R2_INV_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R2_INV_1 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9169));
  sky130_fd_sc_hd__clkbuf_4 T25Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9205));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R0_INV_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9241));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R1_INV_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R2_INV_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R2_INV_1 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9277));
  sky130_fd_sc_hd__clkbuf_4 T25Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9313));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R0_INV_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9349));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R1_INV_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R2_INV_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R2_INV_1 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9385));
  sky130_fd_sc_hd__clkbuf_4 T25Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9421));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R0_INV_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9457));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R1_INV_0 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R2_INV_0 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R2_INV_1 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9493));
  sky130_fd_sc_hd__clkbuf_4 T25Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9529));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R0_INV_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9565));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R1_INV_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R2_INV_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R2_INV_1 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9601));
  sky130_fd_sc_hd__clkbuf_4 T25Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9637));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R0_INV_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9673));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R1_INV_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R2_INV_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R2_INV_1 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9709));
  sky130_fd_sc_hd__clkbuf_4 T25Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B890));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R0_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B926));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R1_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R2_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R2_INV_1 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B962));
  sky130_fd_sc_hd__clkbuf_4 T25Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B998));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R0_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1034));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R1_INV_0 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R2_INV_0 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R2_INV_1 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1070));
  sky130_fd_sc_hd__clkbuf_4 T26Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B36));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R0_INV_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B71));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R1_INV_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R2_INV_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R2_INV_1 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B106));
  sky130_fd_sc_hd__clkbuf_4 T26Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1107));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R0_INV_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1143));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R1_INV_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R2_INV_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R2_INV_1 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1179));
  sky130_fd_sc_hd__clkbuf_4 T26Y11__R0_BUF_0 (.A(clk_L1_B75), .X(clk_L0_B1215));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R0_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1251));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R1_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R2_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R2_INV_1 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1287));
  sky130_fd_sc_hd__clkbuf_4 T26Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1323));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R0_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y12__R1_BUF_0 (.A(clk_L1_B84), .X(clk_L0_B1359));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R1_INV_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R2_INV_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R2_INV_1 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1395));
  sky130_fd_sc_hd__clkbuf_4 T26Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1431));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R0_INV_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1467));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R1_INV_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R2_INV_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R2_INV_1 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y13__R3_BUF_0 (.A(clk_L1_B93), .X(clk_L0_B1503));
  sky130_fd_sc_hd__clkbuf_4 T26Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1539));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R0_INV_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1574));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R1_INV_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R2_INV_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R2_INV_1 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1610));
  sky130_fd_sc_hd__clkbuf_4 T26Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1646));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R0_INV_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1682));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R1_INV_0 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R2_INV_0 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R2_INV_1 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1718));
  sky130_fd_sc_hd__clkbuf_4 T26Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1754));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R0_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1790));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R1_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R2_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R2_INV_1 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1826));
  sky130_fd_sc_hd__clkbuf_4 T26Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1862));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R0_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1898));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R1_INV_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R2_INV_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R2_INV_1 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1934));
  sky130_fd_sc_hd__clkbuf_4 T26Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1970));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R0_INV_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2006));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R1_INV_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R2_INV_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R2_INV_1 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2042));
  sky130_fd_sc_hd__clkbuf_4 T26Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2078));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R0_INV_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2114));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R1_INV_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R2_INV_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R2_INV_1 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2150));
  sky130_fd_sc_hd__clkbuf_4 T26Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B141));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R0_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y1__R1_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B11));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R1_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R2_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R2_INV_1 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B211));
  sky130_fd_sc_hd__clkbuf_4 T26Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2186));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R0_INV_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2222));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R1_INV_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R2_INV_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R2_INV_1 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2258));
  sky130_fd_sc_hd__clkbuf_4 T26Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2294));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R0_INV_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2330));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R1_INV_0 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R2_INV_0 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R2_INV_1 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2366));
  sky130_fd_sc_hd__clkbuf_4 T26Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2402));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R0_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2438));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R1_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R2_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R2_INV_1 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2474));
  sky130_fd_sc_hd__clkbuf_4 T26Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2510));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R0_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2546));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R1_INV_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R2_INV_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R2_INV_1 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2582));
  sky130_fd_sc_hd__clkbuf_4 T26Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2618));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R0_INV_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2654));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R1_INV_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R2_INV_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R2_INV_1 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2690));
  sky130_fd_sc_hd__clkbuf_4 T26Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2726));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R0_INV_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2762));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R1_INV_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R2_INV_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R2_INV_1 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2798));
  sky130_fd_sc_hd__clkbuf_4 T26Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2834));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R0_INV_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2870));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R1_INV_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R2_INV_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R2_INV_1 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2906));
  sky130_fd_sc_hd__clkbuf_4 T26Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2942));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R0_INV_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2978));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R1_INV_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R2_INV_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R2_INV_1 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3014));
  sky130_fd_sc_hd__clkbuf_4 T26Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3050));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R0_INV_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3086));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R1_INV_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R2_INV_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R2_INV_1 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3122));
  sky130_fd_sc_hd__clkbuf_4 T26Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3158));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R0_INV_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3194));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R1_INV_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R2_INV_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R2_INV_1 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3230));
  sky130_fd_sc_hd__clkbuf_4 T26Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B246));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R0_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B281));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R1_INV_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R2_INV_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R2_INV_1 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B317));
  sky130_fd_sc_hd__clkbuf_4 T26Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3266));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R0_INV_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3302));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R1_INV_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R2_INV_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R2_INV_1 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3338));
  sky130_fd_sc_hd__clkbuf_4 T26Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3374));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R0_INV_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3410));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R1_INV_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R2_INV_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R2_INV_1 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3446));
  sky130_fd_sc_hd__clkbuf_4 T26Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3482));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R0_INV_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3518));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R1_INV_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R2_INV_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R2_INV_1 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3554));
  sky130_fd_sc_hd__clkbuf_4 T26Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3590));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R0_INV_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3626));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R1_INV_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R2_INV_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R2_INV_1 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3662));
  sky130_fd_sc_hd__clkbuf_4 T26Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3698));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R0_INV_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3734));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R1_INV_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R2_INV_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R2_INV_1 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3770));
  sky130_fd_sc_hd__clkbuf_4 T26Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3806));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R0_INV_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3842));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R1_INV_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R2_INV_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R2_INV_1 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3878));
  sky130_fd_sc_hd__clkbuf_4 T26Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3914));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R0_INV_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3950));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R1_INV_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R2_INV_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R2_INV_1 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3986));
  sky130_fd_sc_hd__clkbuf_4 T26Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4022));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R0_INV_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4058));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R1_INV_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R2_INV_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R2_INV_1 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4094));
  sky130_fd_sc_hd__clkbuf_4 T26Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4130));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R0_INV_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4166));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R1_INV_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R2_INV_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R2_INV_1 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4202));
  sky130_fd_sc_hd__clkbuf_4 T26Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4238));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R0_INV_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4274));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R1_INV_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R2_INV_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R2_INV_1 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4310));
  sky130_fd_sc_hd__clkbuf_4 T26Y3__R0_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B22));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R0_INV_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B387));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R1_INV_0 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R2_INV_0 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R2_INV_1 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B423));
  sky130_fd_sc_hd__clkbuf_4 T26Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4346));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R0_INV_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4382));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R1_INV_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R2_INV_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R2_INV_1 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4418));
  sky130_fd_sc_hd__clkbuf_4 T26Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4454));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R0_INV_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4490));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R1_INV_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R2_INV_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R2_INV_1 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4526));
  sky130_fd_sc_hd__clkbuf_4 T26Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4562));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R0_INV_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4598));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R1_INV_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R2_INV_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R2_INV_1 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4634));
  sky130_fd_sc_hd__clkbuf_4 T26Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4670));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R0_INV_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4706));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R1_INV_0 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R2_INV_0 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R2_INV_1 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4742));
  sky130_fd_sc_hd__clkbuf_4 T26Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4778));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R0_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4814));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R1_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R2_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R2_INV_1 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4850));
  sky130_fd_sc_hd__clkbuf_4 T26Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4886));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R0_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4922));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R1_INV_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R2_INV_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R2_INV_1 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4958));
  sky130_fd_sc_hd__clkbuf_4 T26Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4994));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R0_INV_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5030));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R1_INV_0 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R2_INV_0 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R2_INV_1 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5066));
  sky130_fd_sc_hd__clkbuf_4 T26Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5102));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R0_INV_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5138));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R1_INV_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R2_INV_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R2_INV_1 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5174));
  sky130_fd_sc_hd__clkbuf_4 T26Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5210));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R0_INV_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5246));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R1_INV_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R2_INV_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R2_INV_1 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5282));
  sky130_fd_sc_hd__clkbuf_4 T26Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5318));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R0_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5354));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R1_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R2_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R2_INV_1 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5390));
  sky130_fd_sc_hd__clkbuf_4 T26Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B459));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R0_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y4__R1_BUF_0 (.A(clk_L1_B30), .X(clk_L0_B495));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R1_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R2_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R2_INV_1 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B531));
  sky130_fd_sc_hd__clkbuf_4 T26Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5426));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R0_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5462));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R1_INV_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R2_INV_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R2_INV_1 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5498));
  sky130_fd_sc_hd__clkbuf_4 T26Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5534));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R0_INV_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5570));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R1_INV_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R2_INV_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R2_INV_1 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5606));
  sky130_fd_sc_hd__clkbuf_4 T26Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5642));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R0_INV_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5678));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R1_INV_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R2_INV_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R2_INV_1 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5714));
  sky130_fd_sc_hd__clkbuf_4 T26Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5750));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R0_INV_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5786));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R1_INV_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R2_INV_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R2_INV_1 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5822));
  sky130_fd_sc_hd__clkbuf_4 T26Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5858));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R0_INV_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5894));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R1_INV_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R2_INV_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R2_INV_1 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5930));
  sky130_fd_sc_hd__clkbuf_4 T26Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5966));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R0_INV_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6002));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R1_INV_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R2_INV_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R2_INV_1 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6038));
  sky130_fd_sc_hd__clkbuf_4 T26Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6074));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R0_INV_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6110));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R1_INV_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R2_INV_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R2_INV_1 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6146));
  sky130_fd_sc_hd__clkbuf_4 T26Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6182));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R0_INV_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6218));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R1_INV_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R2_INV_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R2_INV_1 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6254));
  sky130_fd_sc_hd__clkbuf_4 T26Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6290));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R0_INV_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6326));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R1_INV_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R2_INV_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R2_INV_1 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6362));
  sky130_fd_sc_hd__clkbuf_4 T26Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6398));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R0_INV_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6434));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R1_INV_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R2_INV_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R2_INV_1 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6470));
  sky130_fd_sc_hd__clkbuf_4 T26Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B567));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R0_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B603));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R1_INV_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R2_INV_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R2_INV_1 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y5__R3_BUF_0 (.A(clk_L1_B39), .X(clk_L0_B639));
  sky130_fd_sc_hd__clkbuf_4 T26Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6506));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R0_INV_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6542));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R1_INV_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R2_INV_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R2_INV_1 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6578));
  sky130_fd_sc_hd__clkbuf_4 T26Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6614));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R0_INV_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6650));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R1_INV_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R2_INV_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R2_INV_1 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6686));
  sky130_fd_sc_hd__clkbuf_4 T26Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6722));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R0_INV_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6758));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R1_INV_0 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R2_INV_0 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R2_INV_1 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6794));
  sky130_fd_sc_hd__clkbuf_4 T26Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6830));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R0_INV_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6866));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R1_INV_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R2_INV_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R2_INV_1 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6902));
  sky130_fd_sc_hd__clkbuf_4 T26Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6938));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R0_INV_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6974));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R1_INV_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R2_INV_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R2_INV_1 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7010));
  sky130_fd_sc_hd__clkbuf_4 T26Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7046));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R0_INV_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7082));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R1_INV_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R2_INV_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R2_INV_1 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7118));
  sky130_fd_sc_hd__clkbuf_4 T26Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7154));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R0_INV_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7190));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R1_INV_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R2_INV_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R2_INV_1 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7226));
  sky130_fd_sc_hd__clkbuf_4 T26Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7262));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R0_INV_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7298));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R1_INV_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R2_INV_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R2_INV_1 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7334));
  sky130_fd_sc_hd__clkbuf_4 T26Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7370));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R0_INV_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7406));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R1_INV_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R2_INV_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R2_INV_1 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7442));
  sky130_fd_sc_hd__clkbuf_4 T26Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7478));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R0_INV_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7514));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R1_INV_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R2_INV_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R2_INV_1 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7550));
  sky130_fd_sc_hd__clkbuf_4 T26Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B675));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R0_INV_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B711));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R1_INV_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R2_INV_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R2_INV_1 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B747));
  sky130_fd_sc_hd__clkbuf_4 T26Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7586));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R0_INV_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7622));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R1_INV_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R2_INV_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R2_INV_1 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7658));
  sky130_fd_sc_hd__clkbuf_4 T26Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7694));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R0_INV_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7730));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R1_INV_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R2_INV_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R2_INV_1 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7766));
  sky130_fd_sc_hd__clkbuf_4 T26Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7802));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R0_INV_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7838));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R1_INV_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R2_INV_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R2_INV_1 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7874));
  sky130_fd_sc_hd__clkbuf_4 T26Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7910));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R0_INV_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7946));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R1_INV_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R2_INV_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R2_INV_1 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7982));
  sky130_fd_sc_hd__clkbuf_4 T26Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8018));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R0_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8054));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R1_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R2_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R2_INV_1 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8090));
  sky130_fd_sc_hd__clkbuf_4 T26Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8126));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R0_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8162));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R1_INV_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R2_INV_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R2_INV_1 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8198));
  sky130_fd_sc_hd__clkbuf_4 T26Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8234));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R0_INV_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8270));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R1_INV_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R2_INV_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R2_INV_1 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8306));
  sky130_fd_sc_hd__clkbuf_4 T26Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8342));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R0_INV_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8378));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R1_INV_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R2_INV_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R2_INV_1 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8414));
  sky130_fd_sc_hd__clkbuf_4 T26Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8450));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R0_INV_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8486));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R1_INV_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R2_INV_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R2_INV_1 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8522));
  sky130_fd_sc_hd__clkbuf_4 T26Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8558));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R0_INV_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8594));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R1_INV_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R2_INV_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R2_INV_1 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8630));
  sky130_fd_sc_hd__clkbuf_4 T26Y7__R0_BUF_0 (.A(clk_L1_B48), .X(clk_L0_B783));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R0_INV_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B819));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R1_INV_0 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R2_INV_0 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R2_INV_1 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B855));
  sky130_fd_sc_hd__clkbuf_4 T26Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8666));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R0_INV_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8702));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R1_INV_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R2_INV_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R2_INV_1 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8738));
  sky130_fd_sc_hd__clkbuf_4 T26Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8774));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R0_INV_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8810));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R1_INV_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R2_INV_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R2_INV_1 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8846));
  sky130_fd_sc_hd__clkbuf_4 T26Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8882));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R0_INV_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8918));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R1_INV_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R2_INV_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R2_INV_1 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8954));
  sky130_fd_sc_hd__clkbuf_4 T26Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8990));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R0_INV_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9026));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R1_INV_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R2_INV_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R2_INV_1 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9062));
  sky130_fd_sc_hd__clkbuf_4 T26Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9098));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R0_INV_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9134));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R1_INV_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R2_INV_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R2_INV_1 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9170));
  sky130_fd_sc_hd__clkbuf_4 T26Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9206));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R0_INV_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9242));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R1_INV_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R2_INV_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R2_INV_1 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9278));
  sky130_fd_sc_hd__clkbuf_4 T26Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9314));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R0_INV_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9350));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R1_INV_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R2_INV_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R2_INV_1 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9386));
  sky130_fd_sc_hd__clkbuf_4 T26Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9422));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R0_INV_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9458));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R1_INV_0 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R2_INV_0 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R2_INV_1 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9494));
  sky130_fd_sc_hd__clkbuf_4 T26Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9530));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R0_INV_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9566));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R1_INV_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R2_INV_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R2_INV_1 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9602));
  sky130_fd_sc_hd__clkbuf_4 T26Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9638));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R0_INV_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9674));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R1_INV_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R2_INV_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R2_INV_1 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9710));
  sky130_fd_sc_hd__clkbuf_4 T26Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B891));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R0_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y8__R1_BUF_0 (.A(clk_L1_B57), .X(clk_L0_B927));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R1_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R2_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R2_INV_1 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B963));
  sky130_fd_sc_hd__clkbuf_4 T26Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B999));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R0_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1035));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R1_INV_0 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R2_INV_0 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R2_INV_1 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y9__R3_BUF_0 (.A(clk_L1_B66), .X(clk_L0_B1071));
  sky130_fd_sc_hd__clkbuf_4 T27Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B37));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R0_INV_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B72));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R1_INV_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R2_INV_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R2_INV_1 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B107));
  sky130_fd_sc_hd__clkbuf_4 T27Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1108));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R0_INV_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1144));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R1_INV_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R2_INV_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R2_INV_1 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1180));
  sky130_fd_sc_hd__clkbuf_4 T27Y11__R0_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B76));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R0_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1252));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R1_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R2_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R2_INV_1 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1288));
  sky130_fd_sc_hd__clkbuf_4 T27Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1324));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R0_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y12__R1_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B85));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R1_INV_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R2_INV_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R2_INV_1 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1396));
  sky130_fd_sc_hd__clkbuf_4 T27Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1432));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R0_INV_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1468));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R1_INV_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R2_INV_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R2_INV_1 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y13__R3_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B94));
  sky130_fd_sc_hd__clkbuf_4 T27Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1540));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R0_INV_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1575));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R1_INV_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R2_INV_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R2_INV_1 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1611));
  sky130_fd_sc_hd__clkbuf_4 T27Y15__R0_BUF_0 (.A(clk_L1_B102), .X(clk_L0_B1647));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R0_INV_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1683));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R1_INV_0 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R2_INV_0 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R2_INV_1 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1719));
  sky130_fd_sc_hd__clkbuf_4 T27Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1755));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R0_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y16__R1_BUF_0 (.A(clk_L1_B111), .X(clk_L0_B1791));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R1_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R2_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R2_INV_1 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1827));
  sky130_fd_sc_hd__clkbuf_4 T27Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1863));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R0_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1899));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R1_INV_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R2_INV_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R2_INV_1 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y17__R3_BUF_0 (.A(clk_L1_B120), .X(clk_L0_B1935));
  sky130_fd_sc_hd__clkbuf_4 T27Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1971));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R0_INV_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2007));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R1_INV_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R2_INV_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R2_INV_1 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2043));
  sky130_fd_sc_hd__clkbuf_4 T27Y19__R0_BUF_0 (.A(clk_L1_B129), .X(clk_L0_B2079));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R0_INV_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2115));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R1_INV_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R2_INV_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R2_INV_1 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2151));
  sky130_fd_sc_hd__clkbuf_4 T27Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B142));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R0_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B177));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R1_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R2_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R2_INV_1 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B212));
  sky130_fd_sc_hd__clkbuf_4 T27Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2187));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R0_INV_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y20__R1_BUF_0 (.A(clk_L1_B138), .X(clk_L0_B2223));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R1_INV_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R2_INV_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R2_INV_1 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2259));
  sky130_fd_sc_hd__clkbuf_4 T27Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2295));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R0_INV_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2331));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R1_INV_0 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R2_INV_0 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R2_INV_1 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y21__R3_BUF_0 (.A(clk_L1_B147), .X(clk_L0_B2367));
  sky130_fd_sc_hd__clkbuf_4 T27Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2403));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R0_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2439));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R1_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R2_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R2_INV_1 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2475));
  sky130_fd_sc_hd__clkbuf_4 T27Y23__R0_BUF_0 (.A(clk_L1_B156), .X(clk_L0_B2511));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R0_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2547));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R1_INV_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R2_INV_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R2_INV_1 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2583));
  sky130_fd_sc_hd__clkbuf_4 T27Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2619));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R0_INV_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y24__R1_BUF_0 (.A(clk_L1_B165), .X(clk_L0_B2655));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R1_INV_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R2_INV_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R2_INV_1 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2691));
  sky130_fd_sc_hd__clkbuf_4 T27Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2727));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R0_INV_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2763));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R1_INV_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R2_INV_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R2_INV_1 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y25__R3_BUF_0 (.A(clk_L1_B174), .X(clk_L0_B2799));
  sky130_fd_sc_hd__clkbuf_4 T27Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2835));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R0_INV_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2871));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R1_INV_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R2_INV_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R2_INV_1 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2907));
  sky130_fd_sc_hd__clkbuf_4 T27Y27__R0_BUF_0 (.A(clk_L1_B183), .X(clk_L0_B2943));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R0_INV_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2979));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R1_INV_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R2_INV_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R2_INV_1 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3015));
  sky130_fd_sc_hd__clkbuf_4 T27Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3051));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R0_INV_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y28__R1_BUF_0 (.A(clk_L1_B192), .X(clk_L0_B3087));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R1_INV_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R2_INV_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R2_INV_1 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3123));
  sky130_fd_sc_hd__clkbuf_4 T27Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3159));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R0_INV_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3195));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R1_INV_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R2_INV_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R2_INV_1 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y29__R3_BUF_0 (.A(clk_L1_B201), .X(clk_L0_B3231));
  sky130_fd_sc_hd__clkbuf_4 T27Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B247));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R0_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B282));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R1_INV_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R2_INV_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R2_INV_1 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B318));
  sky130_fd_sc_hd__clkbuf_4 T27Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3267));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R0_INV_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3303));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R1_INV_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R2_INV_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R2_INV_1 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3339));
  sky130_fd_sc_hd__clkbuf_4 T27Y31__R0_BUF_0 (.A(clk_L1_B210), .X(clk_L0_B3375));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R0_INV_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3411));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R1_INV_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R2_INV_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R2_INV_1 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3447));
  sky130_fd_sc_hd__clkbuf_4 T27Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3483));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R0_INV_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y32__R1_BUF_0 (.A(clk_L1_B219), .X(clk_L0_B3519));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R1_INV_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R2_INV_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R2_INV_1 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3555));
  sky130_fd_sc_hd__clkbuf_4 T27Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3591));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R0_INV_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3627));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R1_INV_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R2_INV_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R2_INV_1 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y33__R3_BUF_0 (.A(clk_L1_B228), .X(clk_L0_B3663));
  sky130_fd_sc_hd__clkbuf_4 T27Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3699));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R0_INV_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3735));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R1_INV_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R2_INV_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R2_INV_1 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3771));
  sky130_fd_sc_hd__clkbuf_4 T27Y35__R0_BUF_0 (.A(clk_L1_B237), .X(clk_L0_B3807));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R0_INV_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3843));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R1_INV_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R2_INV_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R2_INV_1 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3879));
  sky130_fd_sc_hd__clkbuf_4 T27Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3915));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R0_INV_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y36__R1_BUF_0 (.A(clk_L1_B246), .X(clk_L0_B3951));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R1_INV_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R2_INV_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R2_INV_1 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3987));
  sky130_fd_sc_hd__clkbuf_4 T27Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4023));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R0_INV_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4059));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R1_INV_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R2_INV_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R2_INV_1 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y37__R3_BUF_0 (.A(clk_L1_B255), .X(clk_L0_B4095));
  sky130_fd_sc_hd__clkbuf_4 T27Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4131));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R0_INV_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4167));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R1_INV_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R2_INV_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R2_INV_1 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4203));
  sky130_fd_sc_hd__clkbuf_4 T27Y39__R0_BUF_0 (.A(clk_L1_B264), .X(clk_L0_B4239));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R0_INV_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4275));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R1_INV_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R2_INV_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R2_INV_1 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4311));
  sky130_fd_sc_hd__clkbuf_4 T27Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B353));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R0_INV_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B388));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R1_INV_0 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R2_INV_0 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R2_INV_1 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B424));
  sky130_fd_sc_hd__clkbuf_4 T27Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4347));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R0_INV_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y40__R1_BUF_0 (.A(clk_L1_B273), .X(clk_L0_B4383));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R1_INV_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R2_INV_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R2_INV_1 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4419));
  sky130_fd_sc_hd__clkbuf_4 T27Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4455));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R0_INV_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4491));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R1_INV_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R2_INV_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R2_INV_1 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y41__R3_BUF_0 (.A(clk_L1_B282), .X(clk_L0_B4527));
  sky130_fd_sc_hd__clkbuf_4 T27Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4563));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R0_INV_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4599));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R1_INV_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R2_INV_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R2_INV_1 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4635));
  sky130_fd_sc_hd__clkbuf_4 T27Y43__R0_BUF_0 (.A(clk_L1_B291), .X(clk_L0_B4671));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R0_INV_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4707));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R1_INV_0 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R2_INV_0 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R2_INV_1 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4743));
  sky130_fd_sc_hd__clkbuf_4 T27Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4779));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R0_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y44__R1_BUF_0 (.A(clk_L1_B300), .X(clk_L0_B4815));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R1_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R2_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R2_INV_1 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4851));
  sky130_fd_sc_hd__clkbuf_4 T27Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4887));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R0_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4923));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R1_INV_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R2_INV_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R2_INV_1 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y45__R3_BUF_0 (.A(clk_L1_B309), .X(clk_L0_B4959));
  sky130_fd_sc_hd__clkbuf_4 T27Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4995));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R0_INV_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5031));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R1_INV_0 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R2_INV_0 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R2_INV_1 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5067));
  sky130_fd_sc_hd__clkbuf_4 T27Y47__R0_BUF_0 (.A(clk_L1_B318), .X(clk_L0_B5103));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R0_INV_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5139));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R1_INV_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R2_INV_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R2_INV_1 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5175));
  sky130_fd_sc_hd__clkbuf_4 T27Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5211));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R0_INV_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y48__R1_BUF_0 (.A(clk_L1_B327), .X(clk_L0_B5247));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R1_INV_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R2_INV_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R2_INV_1 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5283));
  sky130_fd_sc_hd__clkbuf_4 T27Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5319));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R0_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5355));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R1_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R2_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R2_INV_1 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y49__R3_BUF_0 (.A(clk_L1_B336), .X(clk_L0_B5391));
  sky130_fd_sc_hd__clkbuf_4 T27Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B460));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R0_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y4__R1_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B31));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R1_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R2_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R2_INV_1 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B532));
  sky130_fd_sc_hd__clkbuf_4 T27Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5427));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R0_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5463));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R1_INV_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R2_INV_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R2_INV_1 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5499));
  sky130_fd_sc_hd__clkbuf_4 T27Y51__R0_BUF_0 (.A(clk_L1_B345), .X(clk_L0_B5535));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R0_INV_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5571));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R1_INV_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R2_INV_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R2_INV_1 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5607));
  sky130_fd_sc_hd__clkbuf_4 T27Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5643));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R0_INV_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y52__R1_BUF_0 (.A(clk_L1_B354), .X(clk_L0_B5679));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R1_INV_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R2_INV_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R2_INV_1 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5715));
  sky130_fd_sc_hd__clkbuf_4 T27Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5751));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R0_INV_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5787));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R1_INV_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R2_INV_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R2_INV_1 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y53__R3_BUF_0 (.A(clk_L1_B363), .X(clk_L0_B5823));
  sky130_fd_sc_hd__clkbuf_4 T27Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5859));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R0_INV_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5895));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R1_INV_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R2_INV_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R2_INV_1 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5931));
  sky130_fd_sc_hd__clkbuf_4 T27Y55__R0_BUF_0 (.A(clk_L1_B372), .X(clk_L0_B5967));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R0_INV_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6003));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R1_INV_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R2_INV_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R2_INV_1 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6039));
  sky130_fd_sc_hd__clkbuf_4 T27Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6075));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R0_INV_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y56__R1_BUF_0 (.A(clk_L1_B381), .X(clk_L0_B6111));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R1_INV_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R2_INV_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R2_INV_1 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6147));
  sky130_fd_sc_hd__clkbuf_4 T27Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6183));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R0_INV_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6219));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R1_INV_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R2_INV_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R2_INV_1 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y57__R3_BUF_0 (.A(clk_L1_B390), .X(clk_L0_B6255));
  sky130_fd_sc_hd__clkbuf_4 T27Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6291));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R0_INV_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6327));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R1_INV_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R2_INV_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R2_INV_1 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6363));
  sky130_fd_sc_hd__clkbuf_4 T27Y59__R0_BUF_0 (.A(clk_L1_B399), .X(clk_L0_B6399));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R0_INV_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6435));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R1_INV_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R2_INV_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R2_INV_1 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6471));
  sky130_fd_sc_hd__clkbuf_4 T27Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B568));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R0_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B604));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R1_INV_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R2_INV_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R2_INV_1 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y5__R3_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B40));
  sky130_fd_sc_hd__clkbuf_4 T27Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6507));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R0_INV_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y60__R1_BUF_0 (.A(clk_L1_B408), .X(clk_L0_B6543));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R1_INV_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R2_INV_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R2_INV_1 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6579));
  sky130_fd_sc_hd__clkbuf_4 T27Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6615));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R0_INV_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6651));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R1_INV_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R2_INV_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R2_INV_1 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y61__R3_BUF_0 (.A(clk_L1_B417), .X(clk_L0_B6687));
  sky130_fd_sc_hd__clkbuf_4 T27Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6723));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R0_INV_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6759));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R1_INV_0 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R2_INV_0 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R2_INV_1 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6795));
  sky130_fd_sc_hd__clkbuf_4 T27Y63__R0_BUF_0 (.A(clk_L1_B426), .X(clk_L0_B6831));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R0_INV_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6867));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R1_INV_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R2_INV_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R2_INV_1 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6903));
  sky130_fd_sc_hd__clkbuf_4 T27Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6939));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R0_INV_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y64__R1_BUF_0 (.A(clk_L1_B435), .X(clk_L0_B6975));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R1_INV_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R2_INV_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R2_INV_1 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7011));
  sky130_fd_sc_hd__clkbuf_4 T27Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7047));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R0_INV_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7083));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R1_INV_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R2_INV_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R2_INV_1 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y65__R3_BUF_0 (.A(clk_L1_B444), .X(clk_L0_B7119));
  sky130_fd_sc_hd__clkbuf_4 T27Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7155));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R0_INV_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7191));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R1_INV_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R2_INV_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R2_INV_1 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7227));
  sky130_fd_sc_hd__clkbuf_4 T27Y67__R0_BUF_0 (.A(clk_L1_B453), .X(clk_L0_B7263));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R0_INV_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7299));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R1_INV_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R2_INV_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R2_INV_1 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7335));
  sky130_fd_sc_hd__clkbuf_4 T27Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7371));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R0_INV_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y68__R1_BUF_0 (.A(clk_L1_B462), .X(clk_L0_B7407));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R1_INV_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R2_INV_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R2_INV_1 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7443));
  sky130_fd_sc_hd__clkbuf_4 T27Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7479));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R0_INV_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7515));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R1_INV_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R2_INV_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R2_INV_1 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y69__R3_BUF_0 (.A(clk_L1_B471), .X(clk_L0_B7551));
  sky130_fd_sc_hd__clkbuf_4 T27Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B676));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R0_INV_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B712));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R1_INV_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R2_INV_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R2_INV_1 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B748));
  sky130_fd_sc_hd__clkbuf_4 T27Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7587));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R0_INV_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7623));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R1_INV_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R2_INV_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R2_INV_1 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7659));
  sky130_fd_sc_hd__clkbuf_4 T27Y71__R0_BUF_0 (.A(clk_L1_B480), .X(clk_L0_B7695));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R0_INV_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7731));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R1_INV_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R2_INV_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R2_INV_1 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7767));
  sky130_fd_sc_hd__clkbuf_4 T27Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7803));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R0_INV_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y72__R1_BUF_0 (.A(clk_L1_B489), .X(clk_L0_B7839));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R1_INV_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R2_INV_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R2_INV_1 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7875));
  sky130_fd_sc_hd__clkbuf_4 T27Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7911));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R0_INV_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7947));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R1_INV_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R2_INV_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R2_INV_1 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y73__R3_BUF_0 (.A(clk_L1_B498), .X(clk_L0_B7983));
  sky130_fd_sc_hd__clkbuf_4 T27Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8019));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R0_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8055));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R1_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R2_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R2_INV_1 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8091));
  sky130_fd_sc_hd__clkbuf_4 T27Y75__R0_BUF_0 (.A(clk_L1_B507), .X(clk_L0_B8127));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R0_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8163));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R1_INV_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R2_INV_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R2_INV_1 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8199));
  sky130_fd_sc_hd__clkbuf_4 T27Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8235));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R0_INV_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y76__R1_BUF_0 (.A(clk_L1_B516), .X(clk_L0_B8271));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R1_INV_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R2_INV_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R2_INV_1 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8307));
  sky130_fd_sc_hd__clkbuf_4 T27Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8343));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R0_INV_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8379));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R1_INV_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R2_INV_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R2_INV_1 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y77__R3_BUF_0 (.A(clk_L1_B525), .X(clk_L0_B8415));
  sky130_fd_sc_hd__clkbuf_4 T27Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8451));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R0_INV_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8487));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R1_INV_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R2_INV_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R2_INV_1 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8523));
  sky130_fd_sc_hd__clkbuf_4 T27Y79__R0_BUF_0 (.A(clk_L1_B534), .X(clk_L0_B8559));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R0_INV_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8595));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R1_INV_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R2_INV_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R2_INV_1 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8631));
  sky130_fd_sc_hd__clkbuf_4 T27Y7__R0_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B49));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R0_INV_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B820));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R1_INV_0 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R2_INV_0 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R2_INV_1 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B856));
  sky130_fd_sc_hd__clkbuf_4 T27Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8667));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R0_INV_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y80__R1_BUF_0 (.A(clk_L1_B543), .X(clk_L0_B8703));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R1_INV_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R2_INV_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R2_INV_1 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8739));
  sky130_fd_sc_hd__clkbuf_4 T27Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8775));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R0_INV_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8811));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R1_INV_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R2_INV_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R2_INV_1 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y81__R3_BUF_0 (.A(clk_L1_B552), .X(clk_L0_B8847));
  sky130_fd_sc_hd__clkbuf_4 T27Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8883));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R0_INV_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8919));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R1_INV_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R2_INV_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R2_INV_1 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8955));
  sky130_fd_sc_hd__clkbuf_4 T27Y83__R0_BUF_0 (.A(clk_L1_B561), .X(clk_L0_B8991));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R0_INV_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9027));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R1_INV_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R2_INV_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R2_INV_1 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9063));
  sky130_fd_sc_hd__clkbuf_4 T27Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9099));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R0_INV_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y84__R1_BUF_0 (.A(clk_L1_B570), .X(clk_L0_B9135));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R1_INV_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R2_INV_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R2_INV_1 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9171));
  sky130_fd_sc_hd__clkbuf_4 T27Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9207));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R0_INV_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9243));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R1_INV_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R2_INV_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R2_INV_1 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y85__R3_BUF_0 (.A(clk_L1_B579), .X(clk_L0_B9279));
  sky130_fd_sc_hd__clkbuf_4 T27Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9315));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R0_INV_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9351));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R1_INV_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R2_INV_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R2_INV_1 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9387));
  sky130_fd_sc_hd__clkbuf_4 T27Y87__R0_BUF_0 (.A(clk_L1_B588), .X(clk_L0_B9423));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R0_INV_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9459));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R1_INV_0 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R2_INV_0 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R2_INV_1 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9495));
  sky130_fd_sc_hd__clkbuf_4 T27Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9531));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R0_INV_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y88__R1_BUF_0 (.A(clk_L1_B597), .X(clk_L0_B9567));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R1_INV_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R2_INV_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R2_INV_1 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9603));
  sky130_fd_sc_hd__clkbuf_4 T27Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9639));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R0_INV_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9675));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R1_INV_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R2_INV_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R2_INV_1 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y89__R3_BUF_0 (.A(clk_L1_B606), .X(clk_L0_B9711));
  sky130_fd_sc_hd__clkbuf_4 T27Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B892));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R0_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y8__R1_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B58));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R1_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R2_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R2_INV_1 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B964));
  sky130_fd_sc_hd__clkbuf_4 T27Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1000));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R0_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1036));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R1_INV_0 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R2_INV_0 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R2_INV_1 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y9__R3_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B67));
  sky130_fd_sc_hd__clkbuf_4 T28Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B38));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R0_INV_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B73));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R1_INV_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R2_INV_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R2_INV_1 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B108));
  sky130_fd_sc_hd__clkbuf_4 T28Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1109));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R0_INV_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1145));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R1_INV_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R2_INV_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R2_INV_1 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1181));
  sky130_fd_sc_hd__clkbuf_4 T28Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1217));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R0_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1253));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R1_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R2_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R2_INV_1 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1289));
  sky130_fd_sc_hd__clkbuf_4 T28Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1325));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R0_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1361));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R1_INV_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R2_INV_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R2_INV_1 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1397));
  sky130_fd_sc_hd__clkbuf_4 T28Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1433));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R0_INV_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1469));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R1_INV_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R2_INV_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R2_INV_1 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1505));
  sky130_fd_sc_hd__clkbuf_4 T28Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1541));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R0_INV_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1576));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R1_INV_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R2_INV_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R2_INV_1 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1612));
  sky130_fd_sc_hd__clkbuf_4 T28Y15__R0_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B103));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R0_INV_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1684));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R1_INV_0 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R2_INV_0 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R2_INV_1 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1720));
  sky130_fd_sc_hd__clkbuf_4 T28Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1756));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R0_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y16__R1_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B7));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R1_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R2_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R2_INV_1 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1828));
  sky130_fd_sc_hd__clkbuf_4 T28Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1864));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R0_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1900));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R1_INV_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R2_INV_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R2_INV_1 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y17__R3_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B121));
  sky130_fd_sc_hd__clkbuf_4 T28Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1972));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R0_INV_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2008));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R1_INV_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R2_INV_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R2_INV_1 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2044));
  sky130_fd_sc_hd__clkbuf_4 T28Y19__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B130));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R0_INV_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2116));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R1_INV_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R2_INV_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R2_INV_1 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2152));
  sky130_fd_sc_hd__clkbuf_4 T28Y1__R0_BUF_0 (.A(clk_L1_B8), .X(clk_L0_B143));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R0_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B178));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R1_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R2_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R2_INV_1 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B213));
  sky130_fd_sc_hd__clkbuf_4 T28Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2188));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R0_INV_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y20__R1_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B139));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R1_INV_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R2_INV_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R2_INV_1 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2260));
  sky130_fd_sc_hd__clkbuf_4 T28Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2296));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R0_INV_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2332));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R1_INV_0 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R2_INV_0 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R2_INV_1 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y21__R3_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B148));
  sky130_fd_sc_hd__clkbuf_4 T28Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2404));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R0_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2440));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R1_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R2_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R2_INV_1 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2476));
  sky130_fd_sc_hd__clkbuf_4 T28Y23__R0_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B157));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R0_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2548));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R1_INV_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R2_INV_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R2_INV_1 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2584));
  sky130_fd_sc_hd__clkbuf_4 T28Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2620));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R0_INV_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y24__R1_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B166));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R1_INV_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R2_INV_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R2_INV_1 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2692));
  sky130_fd_sc_hd__clkbuf_4 T28Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2728));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R0_INV_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2764));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R1_INV_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R2_INV_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R2_INV_1 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y25__R3_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B175));
  sky130_fd_sc_hd__clkbuf_4 T28Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2836));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R0_INV_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2872));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R1_INV_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R2_INV_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R2_INV_1 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2908));
  sky130_fd_sc_hd__clkbuf_4 T28Y27__R0_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B184));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R0_INV_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2980));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R1_INV_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R2_INV_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R2_INV_1 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3016));
  sky130_fd_sc_hd__clkbuf_4 T28Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3052));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R0_INV_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y28__R1_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B193));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R1_INV_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R2_INV_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R2_INV_1 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3124));
  sky130_fd_sc_hd__clkbuf_4 T28Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3160));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R0_INV_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3196));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R1_INV_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R2_INV_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R2_INV_1 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y29__R3_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B202));
  sky130_fd_sc_hd__clkbuf_4 T28Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B248));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R0_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B283));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R1_INV_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R2_INV_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R2_INV_1 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y2__R3_BUF_0 (.A(clk_L1_B19), .X(clk_L0_B319));
  sky130_fd_sc_hd__clkbuf_4 T28Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3268));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R0_INV_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3304));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R1_INV_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R2_INV_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R2_INV_1 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3340));
  sky130_fd_sc_hd__clkbuf_4 T28Y31__R0_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B211));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R0_INV_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3412));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R1_INV_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R2_INV_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R2_INV_1 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3448));
  sky130_fd_sc_hd__clkbuf_4 T28Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3484));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R0_INV_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y32__R1_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B220));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R1_INV_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R2_INV_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R2_INV_1 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3556));
  sky130_fd_sc_hd__clkbuf_4 T28Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3592));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R0_INV_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3628));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R1_INV_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R2_INV_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R2_INV_1 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y33__R3_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B229));
  sky130_fd_sc_hd__clkbuf_4 T28Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3700));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R0_INV_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3736));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R1_INV_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R2_INV_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R2_INV_1 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3772));
  sky130_fd_sc_hd__clkbuf_4 T28Y35__R0_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B238));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R0_INV_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3844));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R1_INV_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R2_INV_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R2_INV_1 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3880));
  sky130_fd_sc_hd__clkbuf_4 T28Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3916));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R0_INV_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y36__R1_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B247));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R1_INV_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R2_INV_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R2_INV_1 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3988));
  sky130_fd_sc_hd__clkbuf_4 T28Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4024));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R0_INV_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4060));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R1_INV_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R2_INV_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R2_INV_1 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y37__R3_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B16));
  sky130_fd_sc_hd__clkbuf_4 T28Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4132));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R0_INV_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4168));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R1_INV_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R2_INV_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R2_INV_1 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4204));
  sky130_fd_sc_hd__clkbuf_4 T28Y39__R0_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B265));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R0_INV_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4276));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R1_INV_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R2_INV_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R2_INV_1 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4312));
  sky130_fd_sc_hd__clkbuf_4 T28Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B354));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R0_INV_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B389));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R1_INV_0 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R2_INV_0 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R2_INV_1 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B425));
  sky130_fd_sc_hd__clkbuf_4 T28Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4348));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R0_INV_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y40__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B274));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R1_INV_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R2_INV_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R2_INV_1 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4420));
  sky130_fd_sc_hd__clkbuf_4 T28Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4456));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R0_INV_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4492));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R1_INV_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R2_INV_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R2_INV_1 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y41__R3_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B283));
  sky130_fd_sc_hd__clkbuf_4 T28Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4564));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R0_INV_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4600));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R1_INV_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R2_INV_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R2_INV_1 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4636));
  sky130_fd_sc_hd__clkbuf_4 T28Y43__R0_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B292));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R0_INV_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4708));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R1_INV_0 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R2_INV_0 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R2_INV_1 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4744));
  sky130_fd_sc_hd__clkbuf_4 T28Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4780));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R0_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y44__R1_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B301));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R1_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R2_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R2_INV_1 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4852));
  sky130_fd_sc_hd__clkbuf_4 T28Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4888));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R0_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4924));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R1_INV_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R2_INV_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R2_INV_1 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y45__R3_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B310));
  sky130_fd_sc_hd__clkbuf_4 T28Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4996));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R0_INV_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5032));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R1_INV_0 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R2_INV_0 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R2_INV_1 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5068));
  sky130_fd_sc_hd__clkbuf_4 T28Y47__R0_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B319));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R0_INV_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5140));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R1_INV_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R2_INV_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R2_INV_1 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5176));
  sky130_fd_sc_hd__clkbuf_4 T28Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5212));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R0_INV_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y48__R1_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B328));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R1_INV_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R2_INV_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R2_INV_1 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5284));
  sky130_fd_sc_hd__clkbuf_4 T28Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5320));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R0_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5356));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R1_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R2_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R2_INV_1 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y49__R3_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B337));
  sky130_fd_sc_hd__clkbuf_4 T28Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B461));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R0_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B497));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R1_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R2_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R2_INV_1 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B533));
  sky130_fd_sc_hd__clkbuf_4 T28Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5428));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R0_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5464));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R1_INV_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R2_INV_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R2_INV_1 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5500));
  sky130_fd_sc_hd__clkbuf_4 T28Y51__R0_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B346));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R0_INV_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5572));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R1_INV_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R2_INV_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R2_INV_1 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5608));
  sky130_fd_sc_hd__clkbuf_4 T28Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5644));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R0_INV_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y52__R1_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B355));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R1_INV_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R2_INV_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R2_INV_1 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5716));
  sky130_fd_sc_hd__clkbuf_4 T28Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5752));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R0_INV_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5788));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R1_INV_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R2_INV_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R2_INV_1 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y53__R3_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B364));
  sky130_fd_sc_hd__clkbuf_4 T28Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5860));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R0_INV_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5896));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R1_INV_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R2_INV_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R2_INV_1 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5932));
  sky130_fd_sc_hd__clkbuf_4 T28Y55__R0_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B373));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R0_INV_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6004));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R1_INV_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R2_INV_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R2_INV_1 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6040));
  sky130_fd_sc_hd__clkbuf_4 T28Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6076));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R0_INV_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y56__R1_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B382));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R1_INV_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R2_INV_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R2_INV_1 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6148));
  sky130_fd_sc_hd__clkbuf_4 T28Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6184));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R0_INV_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6220));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R1_INV_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R2_INV_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R2_INV_1 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y57__R3_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B391));
  sky130_fd_sc_hd__clkbuf_4 T28Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6292));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R0_INV_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6328));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R1_INV_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R2_INV_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R2_INV_1 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6364));
  sky130_fd_sc_hd__clkbuf_4 T28Y59__R0_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B25));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R0_INV_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6436));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R1_INV_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R2_INV_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R2_INV_1 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6472));
  sky130_fd_sc_hd__clkbuf_4 T28Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B569));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R0_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B605));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R1_INV_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R2_INV_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R2_INV_1 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B641));
  sky130_fd_sc_hd__clkbuf_4 T28Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6508));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R0_INV_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y60__R1_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B409));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R1_INV_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R2_INV_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R2_INV_1 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6580));
  sky130_fd_sc_hd__clkbuf_4 T28Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6616));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R0_INV_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6652));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R1_INV_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R2_INV_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R2_INV_1 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y61__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B418));
  sky130_fd_sc_hd__clkbuf_4 T28Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6724));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R0_INV_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6760));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R1_INV_0 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R2_INV_0 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R2_INV_1 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6796));
  sky130_fd_sc_hd__clkbuf_4 T28Y63__R0_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B427));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R0_INV_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6868));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R1_INV_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R2_INV_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R2_INV_1 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6904));
  sky130_fd_sc_hd__clkbuf_4 T28Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6940));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R0_INV_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y64__R1_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B436));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R1_INV_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R2_INV_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R2_INV_1 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7012));
  sky130_fd_sc_hd__clkbuf_4 T28Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7048));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R0_INV_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7084));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R1_INV_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R2_INV_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R2_INV_1 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y65__R3_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B445));
  sky130_fd_sc_hd__clkbuf_4 T28Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7156));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R0_INV_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7192));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R1_INV_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R2_INV_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R2_INV_1 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7228));
  sky130_fd_sc_hd__clkbuf_4 T28Y67__R0_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B454));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R0_INV_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7300));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R1_INV_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R2_INV_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R2_INV_1 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7336));
  sky130_fd_sc_hd__clkbuf_4 T28Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7372));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R0_INV_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y68__R1_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B463));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R1_INV_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R2_INV_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R2_INV_1 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7444));
  sky130_fd_sc_hd__clkbuf_4 T28Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7480));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R0_INV_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7516));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R1_INV_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R2_INV_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R2_INV_1 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y69__R3_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B472));
  sky130_fd_sc_hd__clkbuf_4 T28Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B677));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R0_INV_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B713));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R1_INV_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R2_INV_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R2_INV_1 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B749));
  sky130_fd_sc_hd__clkbuf_4 T28Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7588));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R0_INV_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7624));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R1_INV_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R2_INV_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R2_INV_1 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7660));
  sky130_fd_sc_hd__clkbuf_4 T28Y71__R0_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B481));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R0_INV_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7732));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R1_INV_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R2_INV_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R2_INV_1 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7768));
  sky130_fd_sc_hd__clkbuf_4 T28Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7804));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R0_INV_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y72__R1_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B490));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R1_INV_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R2_INV_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R2_INV_1 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7876));
  sky130_fd_sc_hd__clkbuf_4 T28Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7912));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R0_INV_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7948));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R1_INV_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R2_INV_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R2_INV_1 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y73__R3_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B499));
  sky130_fd_sc_hd__clkbuf_4 T28Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8020));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R0_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8056));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R1_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R2_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R2_INV_1 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8092));
  sky130_fd_sc_hd__clkbuf_4 T28Y75__R0_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B508));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R0_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8164));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R1_INV_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R2_INV_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R2_INV_1 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8200));
  sky130_fd_sc_hd__clkbuf_4 T28Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8236));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R0_INV_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y76__R1_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B517));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R1_INV_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R2_INV_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R2_INV_1 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8308));
  sky130_fd_sc_hd__clkbuf_4 T28Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8344));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R0_INV_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8380));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R1_INV_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R2_INV_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R2_INV_1 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y77__R3_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B526));
  sky130_fd_sc_hd__clkbuf_4 T28Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8452));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R0_INV_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8488));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R1_INV_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R2_INV_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R2_INV_1 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8524));
  sky130_fd_sc_hd__clkbuf_4 T28Y79__R0_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B535));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R0_INV_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8596));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R1_INV_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R2_INV_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R2_INV_1 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8632));
  sky130_fd_sc_hd__clkbuf_4 T28Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B785));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R0_INV_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B821));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R1_INV_0 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R2_INV_0 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R2_INV_1 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B857));
  sky130_fd_sc_hd__clkbuf_4 T28Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8668));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R0_INV_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y80__R1_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B34));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R1_INV_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R2_INV_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R2_INV_1 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8740));
  sky130_fd_sc_hd__clkbuf_4 T28Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8776));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R0_INV_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8812));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R1_INV_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R2_INV_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R2_INV_1 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y81__R3_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B553));
  sky130_fd_sc_hd__clkbuf_4 T28Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8884));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R0_INV_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8920));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R1_INV_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R2_INV_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R2_INV_1 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8956));
  sky130_fd_sc_hd__clkbuf_4 T28Y83__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B562));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R0_INV_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9028));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R1_INV_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R2_INV_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R2_INV_1 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9064));
  sky130_fd_sc_hd__clkbuf_4 T28Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9100));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R0_INV_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y84__R1_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B571));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R1_INV_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R2_INV_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R2_INV_1 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9172));
  sky130_fd_sc_hd__clkbuf_4 T28Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9208));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R0_INV_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9244));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R1_INV_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R2_INV_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R2_INV_1 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y85__R3_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B580));
  sky130_fd_sc_hd__clkbuf_4 T28Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9316));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R0_INV_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9352));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R1_INV_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R2_INV_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R2_INV_1 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9388));
  sky130_fd_sc_hd__clkbuf_4 T28Y87__R0_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B589));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R0_INV_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9460));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R1_INV_0 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R2_INV_0 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R2_INV_1 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9496));
  sky130_fd_sc_hd__clkbuf_4 T28Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9532));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R0_INV_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y88__R1_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B598));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R1_INV_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R2_INV_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R2_INV_1 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9604));
  sky130_fd_sc_hd__clkbuf_4 T28Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9640));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R0_INV_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9676));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R1_INV_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R2_INV_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R2_INV_1 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y89__R3_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B607));
  sky130_fd_sc_hd__clkbuf_4 T28Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B893));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R0_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B929));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R1_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R2_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R2_INV_1 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B965));
  sky130_fd_sc_hd__clkbuf_4 T28Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1001));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R0_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1037));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R1_INV_0 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R2_INV_0 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R2_INV_1 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1073));
  sky130_fd_sc_hd__clkbuf_4 T29Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B39));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R0_INV_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B74));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R1_INV_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R2_INV_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R2_INV_1 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B109));
  sky130_fd_sc_hd__clkbuf_4 T29Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1110));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R0_INV_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1146));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R1_INV_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R2_INV_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R2_INV_1 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1182));
  sky130_fd_sc_hd__clkbuf_4 T29Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1218));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R0_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1254));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R1_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R2_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R2_INV_1 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1290));
  sky130_fd_sc_hd__clkbuf_4 T29Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1326));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R0_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1362));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R1_INV_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R2_INV_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R2_INV_1 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1398));
  sky130_fd_sc_hd__clkbuf_4 T29Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1434));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R0_INV_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1470));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R1_INV_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R2_INV_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R2_INV_1 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1506));
  sky130_fd_sc_hd__clkbuf_4 T29Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1542));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R0_INV_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1577));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R1_INV_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R2_INV_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R2_INV_1 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1613));
  sky130_fd_sc_hd__clkbuf_4 T29Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1649));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R0_INV_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1685));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R1_INV_0 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R2_INV_0 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R2_INV_1 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1721));
  sky130_fd_sc_hd__clkbuf_4 T29Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1757));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R0_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1793));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R1_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R2_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R2_INV_1 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1829));
  sky130_fd_sc_hd__clkbuf_4 T29Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1865));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R0_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1901));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R1_INV_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R2_INV_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R2_INV_1 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1937));
  sky130_fd_sc_hd__clkbuf_4 T29Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1973));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R0_INV_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2009));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R1_INV_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R2_INV_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R2_INV_1 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2045));
  sky130_fd_sc_hd__clkbuf_4 T29Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2081));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R0_INV_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2117));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R1_INV_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R2_INV_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R2_INV_1 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2153));
  sky130_fd_sc_hd__clkbuf_4 T29Y1__R0_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B9));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R0_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B179));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R1_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R2_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R2_INV_1 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B214));
  sky130_fd_sc_hd__clkbuf_4 T29Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2189));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R0_INV_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2225));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R1_INV_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R2_INV_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R2_INV_1 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2261));
  sky130_fd_sc_hd__clkbuf_4 T29Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2297));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R0_INV_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2333));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R1_INV_0 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R2_INV_0 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R2_INV_1 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2369));
  sky130_fd_sc_hd__clkbuf_4 T29Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2405));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R0_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2441));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R1_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R2_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R2_INV_1 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2477));
  sky130_fd_sc_hd__clkbuf_4 T29Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2513));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R0_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2549));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R1_INV_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R2_INV_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R2_INV_1 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2585));
  sky130_fd_sc_hd__clkbuf_4 T29Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2621));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R0_INV_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2657));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R1_INV_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R2_INV_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R2_INV_1 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2693));
  sky130_fd_sc_hd__clkbuf_4 T29Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2729));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R0_INV_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2765));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R1_INV_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R2_INV_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R2_INV_1 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2801));
  sky130_fd_sc_hd__clkbuf_4 T29Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2837));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R0_INV_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2873));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R1_INV_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R2_INV_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R2_INV_1 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2909));
  sky130_fd_sc_hd__clkbuf_4 T29Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2945));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R0_INV_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2981));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R1_INV_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R2_INV_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R2_INV_1 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3017));
  sky130_fd_sc_hd__clkbuf_4 T29Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3053));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R0_INV_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3089));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R1_INV_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R2_INV_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R2_INV_1 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3125));
  sky130_fd_sc_hd__clkbuf_4 T29Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3161));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R0_INV_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3197));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R1_INV_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R2_INV_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R2_INV_1 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3233));
  sky130_fd_sc_hd__clkbuf_4 T29Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B249));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R0_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B284));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R1_INV_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R2_INV_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R2_INV_1 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y2__R3_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B20));
  sky130_fd_sc_hd__clkbuf_4 T29Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3269));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R0_INV_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3305));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R1_INV_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R2_INV_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R2_INV_1 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3341));
  sky130_fd_sc_hd__clkbuf_4 T29Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3377));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R0_INV_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3413));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R1_INV_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R2_INV_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R2_INV_1 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3449));
  sky130_fd_sc_hd__clkbuf_4 T29Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3485));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R0_INV_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3521));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R1_INV_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R2_INV_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R2_INV_1 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3557));
  sky130_fd_sc_hd__clkbuf_4 T29Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3593));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R0_INV_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3629));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R1_INV_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R2_INV_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R2_INV_1 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3665));
  sky130_fd_sc_hd__clkbuf_4 T29Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3701));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R0_INV_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3737));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R1_INV_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R2_INV_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R2_INV_1 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3773));
  sky130_fd_sc_hd__clkbuf_4 T29Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3809));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R0_INV_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3845));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R1_INV_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R2_INV_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R2_INV_1 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3881));
  sky130_fd_sc_hd__clkbuf_4 T29Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3917));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R0_INV_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3953));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R1_INV_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R2_INV_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R2_INV_1 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3989));
  sky130_fd_sc_hd__clkbuf_4 T29Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4025));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R0_INV_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4061));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R1_INV_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R2_INV_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R2_INV_1 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4097));
  sky130_fd_sc_hd__clkbuf_4 T29Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4133));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R0_INV_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4169));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R1_INV_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R2_INV_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R2_INV_1 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4205));
  sky130_fd_sc_hd__clkbuf_4 T29Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4241));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R0_INV_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4277));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R1_INV_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R2_INV_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R2_INV_1 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4313));
  sky130_fd_sc_hd__clkbuf_4 T29Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B355));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R0_INV_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B390));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R1_INV_0 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R2_INV_0 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R2_INV_1 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B426));
  sky130_fd_sc_hd__clkbuf_4 T29Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4349));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R0_INV_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4385));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R1_INV_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R2_INV_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R2_INV_1 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4421));
  sky130_fd_sc_hd__clkbuf_4 T29Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4457));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R0_INV_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4493));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R1_INV_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R2_INV_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R2_INV_1 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4529));
  sky130_fd_sc_hd__clkbuf_4 T29Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4565));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R0_INV_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4601));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R1_INV_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R2_INV_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R2_INV_1 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4637));
  sky130_fd_sc_hd__clkbuf_4 T29Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4673));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R0_INV_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4709));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R1_INV_0 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R2_INV_0 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R2_INV_1 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4745));
  sky130_fd_sc_hd__clkbuf_4 T29Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4781));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R0_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4817));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R1_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R2_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R2_INV_1 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4853));
  sky130_fd_sc_hd__clkbuf_4 T29Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4889));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R0_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4925));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R1_INV_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R2_INV_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R2_INV_1 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4961));
  sky130_fd_sc_hd__clkbuf_4 T29Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4997));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R0_INV_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5033));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R1_INV_0 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R2_INV_0 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R2_INV_1 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5069));
  sky130_fd_sc_hd__clkbuf_4 T29Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5105));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R0_INV_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5141));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R1_INV_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R2_INV_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R2_INV_1 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5177));
  sky130_fd_sc_hd__clkbuf_4 T29Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5213));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R0_INV_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5249));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R1_INV_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R2_INV_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R2_INV_1 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5285));
  sky130_fd_sc_hd__clkbuf_4 T29Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5321));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R0_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5357));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R1_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R2_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R2_INV_1 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5393));
  sky130_fd_sc_hd__clkbuf_4 T29Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B462));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R0_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B498));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R1_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R2_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R2_INV_1 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B534));
  sky130_fd_sc_hd__clkbuf_4 T29Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5429));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R0_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5465));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R1_INV_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R2_INV_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R2_INV_1 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5501));
  sky130_fd_sc_hd__clkbuf_4 T29Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5537));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R0_INV_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5573));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R1_INV_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R2_INV_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R2_INV_1 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5609));
  sky130_fd_sc_hd__clkbuf_4 T29Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5645));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R0_INV_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5681));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R1_INV_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R2_INV_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R2_INV_1 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5717));
  sky130_fd_sc_hd__clkbuf_4 T29Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5753));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R0_INV_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5789));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R1_INV_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R2_INV_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R2_INV_1 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5825));
  sky130_fd_sc_hd__clkbuf_4 T29Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5861));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R0_INV_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5897));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R1_INV_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R2_INV_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R2_INV_1 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5933));
  sky130_fd_sc_hd__clkbuf_4 T29Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5969));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R0_INV_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6005));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R1_INV_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R2_INV_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R2_INV_1 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6041));
  sky130_fd_sc_hd__clkbuf_4 T29Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6077));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R0_INV_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6113));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R1_INV_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R2_INV_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R2_INV_1 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6149));
  sky130_fd_sc_hd__clkbuf_4 T29Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6185));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R0_INV_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6221));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R1_INV_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R2_INV_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R2_INV_1 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6257));
  sky130_fd_sc_hd__clkbuf_4 T29Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6293));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R0_INV_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6329));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R1_INV_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R2_INV_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R2_INV_1 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6365));
  sky130_fd_sc_hd__clkbuf_4 T29Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6401));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R0_INV_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6437));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R1_INV_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R2_INV_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R2_INV_1 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6473));
  sky130_fd_sc_hd__clkbuf_4 T29Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B570));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R0_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B606));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R1_INV_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R2_INV_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R2_INV_1 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B642));
  sky130_fd_sc_hd__clkbuf_4 T29Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6509));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R0_INV_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6545));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R1_INV_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R2_INV_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R2_INV_1 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6581));
  sky130_fd_sc_hd__clkbuf_4 T29Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6617));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R0_INV_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6653));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R1_INV_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R2_INV_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R2_INV_1 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6689));
  sky130_fd_sc_hd__clkbuf_4 T29Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6725));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R0_INV_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6761));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R1_INV_0 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R2_INV_0 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R2_INV_1 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6797));
  sky130_fd_sc_hd__clkbuf_4 T29Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6833));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R0_INV_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6869));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R1_INV_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R2_INV_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R2_INV_1 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6905));
  sky130_fd_sc_hd__clkbuf_4 T29Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6941));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R0_INV_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6977));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R1_INV_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R2_INV_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R2_INV_1 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7013));
  sky130_fd_sc_hd__clkbuf_4 T29Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7049));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R0_INV_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7085));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R1_INV_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R2_INV_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R2_INV_1 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7121));
  sky130_fd_sc_hd__clkbuf_4 T29Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7157));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R0_INV_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7193));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R1_INV_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R2_INV_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R2_INV_1 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7229));
  sky130_fd_sc_hd__clkbuf_4 T29Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7265));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R0_INV_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7301));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R1_INV_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R2_INV_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R2_INV_1 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7337));
  sky130_fd_sc_hd__clkbuf_4 T29Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7373));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R0_INV_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7409));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R1_INV_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R2_INV_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R2_INV_1 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7445));
  sky130_fd_sc_hd__clkbuf_4 T29Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7481));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R0_INV_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7517));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R1_INV_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R2_INV_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R2_INV_1 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7553));
  sky130_fd_sc_hd__clkbuf_4 T29Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B678));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R0_INV_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B714));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R1_INV_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R2_INV_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R2_INV_1 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B750));
  sky130_fd_sc_hd__clkbuf_4 T29Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7589));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R0_INV_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7625));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R1_INV_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R2_INV_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R2_INV_1 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7661));
  sky130_fd_sc_hd__clkbuf_4 T29Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7697));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R0_INV_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7733));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R1_INV_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R2_INV_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R2_INV_1 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7769));
  sky130_fd_sc_hd__clkbuf_4 T29Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7805));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R0_INV_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7841));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R1_INV_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R2_INV_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R2_INV_1 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7877));
  sky130_fd_sc_hd__clkbuf_4 T29Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7913));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R0_INV_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7949));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R1_INV_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R2_INV_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R2_INV_1 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7985));
  sky130_fd_sc_hd__clkbuf_4 T29Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8021));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R0_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8057));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R1_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R2_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R2_INV_1 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8093));
  sky130_fd_sc_hd__clkbuf_4 T29Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8129));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R0_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8165));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R1_INV_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R2_INV_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R2_INV_1 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8201));
  sky130_fd_sc_hd__clkbuf_4 T29Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8237));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R0_INV_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8273));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R1_INV_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R2_INV_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R2_INV_1 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8309));
  sky130_fd_sc_hd__clkbuf_4 T29Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8345));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R0_INV_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8381));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R1_INV_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R2_INV_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R2_INV_1 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8417));
  sky130_fd_sc_hd__clkbuf_4 T29Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8453));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R0_INV_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8489));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R1_INV_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R2_INV_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R2_INV_1 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8525));
  sky130_fd_sc_hd__clkbuf_4 T29Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8561));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R0_INV_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8597));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R1_INV_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R2_INV_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R2_INV_1 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8633));
  sky130_fd_sc_hd__clkbuf_4 T29Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B786));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R0_INV_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B822));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R1_INV_0 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R2_INV_0 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R2_INV_1 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B858));
  sky130_fd_sc_hd__clkbuf_4 T29Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8669));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R0_INV_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8705));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R1_INV_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R2_INV_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R2_INV_1 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8741));
  sky130_fd_sc_hd__clkbuf_4 T29Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8777));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R0_INV_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8813));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R1_INV_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R2_INV_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R2_INV_1 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8849));
  sky130_fd_sc_hd__clkbuf_4 T29Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8885));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R0_INV_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8921));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R1_INV_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R2_INV_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R2_INV_1 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8957));
  sky130_fd_sc_hd__clkbuf_4 T29Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8993));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R0_INV_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9029));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R1_INV_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R2_INV_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R2_INV_1 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9065));
  sky130_fd_sc_hd__clkbuf_4 T29Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9101));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R0_INV_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9137));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R1_INV_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R2_INV_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R2_INV_1 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9173));
  sky130_fd_sc_hd__clkbuf_4 T29Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9209));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R0_INV_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9245));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R1_INV_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R2_INV_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R2_INV_1 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9281));
  sky130_fd_sc_hd__clkbuf_4 T29Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9317));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R0_INV_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9353));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R1_INV_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R2_INV_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R2_INV_1 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9389));
  sky130_fd_sc_hd__clkbuf_4 T29Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9425));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R0_INV_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9461));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R1_INV_0 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R2_INV_0 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R2_INV_1 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9497));
  sky130_fd_sc_hd__clkbuf_4 T29Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9533));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R0_INV_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9569));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R1_INV_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R2_INV_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R2_INV_1 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9605));
  sky130_fd_sc_hd__clkbuf_4 T29Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9641));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R0_INV_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9677));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R1_INV_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R2_INV_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R2_INV_1 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9713));
  sky130_fd_sc_hd__clkbuf_4 T29Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B894));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R0_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B930));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R1_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R2_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R2_INV_1 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B966));
  sky130_fd_sc_hd__clkbuf_4 T29Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1002));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R0_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1038));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R1_INV_0 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R2_INV_0 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R2_INV_1 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1074));
  sky130_fd_sc_hd__clkbuf_4 T2Y0__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B12));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R0_INV_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y0__R1_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B47));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R1_INV_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R2_INV_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R2_INV_1 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B82));
  sky130_fd_sc_hd__clkbuf_4 T2Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1083));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R0_INV_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y10__R1_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1119));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R1_INV_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R2_INV_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R2_INV_1 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1155));
  sky130_fd_sc_hd__clkbuf_4 T2Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1191));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R0_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1227));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R1_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R2_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R2_INV_1 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y11__R3_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1263));
  sky130_fd_sc_hd__clkbuf_4 T2Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1299));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R0_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1335));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R1_INV_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R2_INV_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R2_INV_1 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1371));
  sky130_fd_sc_hd__clkbuf_4 T2Y13__R0_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1407));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R0_INV_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1443));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R1_INV_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R2_INV_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R2_INV_1 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1479));
  sky130_fd_sc_hd__clkbuf_4 T2Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1515));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R0_INV_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y14__R1_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1550));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R1_INV_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R2_INV_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R2_INV_1 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1586));
  sky130_fd_sc_hd__clkbuf_4 T2Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1622));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R0_INV_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1658));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R1_INV_0 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R2_INV_0 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R2_INV_1 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y15__R3_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1694));
  sky130_fd_sc_hd__clkbuf_4 T2Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1730));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R0_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1766));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R1_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R2_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R2_INV_1 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1802));
  sky130_fd_sc_hd__clkbuf_4 T2Y17__R0_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1838));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R0_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1874));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R1_INV_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R2_INV_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R2_INV_1 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1910));
  sky130_fd_sc_hd__clkbuf_4 T2Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1946));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R0_INV_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y18__R1_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1982));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R1_INV_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R2_INV_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R2_INV_1 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2018));
  sky130_fd_sc_hd__clkbuf_4 T2Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2054));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R0_INV_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2090));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R1_INV_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R2_INV_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R2_INV_1 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y19__R3_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2126));
  sky130_fd_sc_hd__clkbuf_4 T2Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B117));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R0_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B152));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R1_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R2_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R2_INV_1 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B187));
  sky130_fd_sc_hd__clkbuf_4 T2Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2162));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R0_INV_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2198));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R1_INV_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R2_INV_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R2_INV_1 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2234));
  sky130_fd_sc_hd__clkbuf_4 T2Y21__R0_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2270));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R0_INV_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2306));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R1_INV_0 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R2_INV_0 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R2_INV_1 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2342));
  sky130_fd_sc_hd__clkbuf_4 T2Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2378));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R0_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y22__R1_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2414));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R1_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R2_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R2_INV_1 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2450));
  sky130_fd_sc_hd__clkbuf_4 T2Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2486));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R0_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2522));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R1_INV_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R2_INV_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R2_INV_1 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y23__R3_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2558));
  sky130_fd_sc_hd__clkbuf_4 T2Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2594));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R0_INV_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2630));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R1_INV_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R2_INV_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R2_INV_1 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2666));
  sky130_fd_sc_hd__clkbuf_4 T2Y25__R0_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2702));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R0_INV_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2738));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R1_INV_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R2_INV_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R2_INV_1 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2774));
  sky130_fd_sc_hd__clkbuf_4 T2Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2810));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R0_INV_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y26__R1_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2846));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R1_INV_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R2_INV_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R2_INV_1 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2882));
  sky130_fd_sc_hd__clkbuf_4 T2Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2918));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R0_INV_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2954));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R1_INV_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R2_INV_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R2_INV_1 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y27__R3_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2990));
  sky130_fd_sc_hd__clkbuf_4 T2Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3026));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R0_INV_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3062));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R1_INV_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R2_INV_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R2_INV_1 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3098));
  sky130_fd_sc_hd__clkbuf_4 T2Y29__R0_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3134));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R0_INV_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3170));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R1_INV_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R2_INV_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R2_INV_1 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3206));
  sky130_fd_sc_hd__clkbuf_4 T2Y2__R0_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B222));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R0_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B257));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R1_INV_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R2_INV_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R2_INV_1 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B293));
  sky130_fd_sc_hd__clkbuf_4 T2Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3242));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R0_INV_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y30__R1_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3278));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R1_INV_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R2_INV_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R2_INV_1 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3314));
  sky130_fd_sc_hd__clkbuf_4 T2Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3350));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R0_INV_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3386));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R1_INV_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R2_INV_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R2_INV_1 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y31__R3_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3422));
  sky130_fd_sc_hd__clkbuf_4 T2Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3458));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R0_INV_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3494));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R1_INV_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R2_INV_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R2_INV_1 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3530));
  sky130_fd_sc_hd__clkbuf_4 T2Y33__R0_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3566));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R0_INV_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3602));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R1_INV_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R2_INV_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R2_INV_1 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3638));
  sky130_fd_sc_hd__clkbuf_4 T2Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3674));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R0_INV_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y34__R1_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3710));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R1_INV_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R2_INV_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R2_INV_1 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3746));
  sky130_fd_sc_hd__clkbuf_4 T2Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3782));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R0_INV_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3818));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R1_INV_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R2_INV_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R2_INV_1 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y35__R3_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3854));
  sky130_fd_sc_hd__clkbuf_4 T2Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3890));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R0_INV_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3926));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R1_INV_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R2_INV_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R2_INV_1 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3962));
  sky130_fd_sc_hd__clkbuf_4 T2Y37__R0_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3998));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R0_INV_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4034));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R1_INV_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R2_INV_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R2_INV_1 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4070));
  sky130_fd_sc_hd__clkbuf_4 T2Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4106));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R0_INV_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y38__R1_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4142));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R1_INV_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R2_INV_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R2_INV_1 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4178));
  sky130_fd_sc_hd__clkbuf_4 T2Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4214));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R0_INV_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4250));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R1_INV_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R2_INV_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R2_INV_1 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y39__R3_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4286));
  sky130_fd_sc_hd__clkbuf_4 T2Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B328));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R0_INV_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B363));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R1_INV_0 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R2_INV_0 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R2_INV_1 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y3__R3_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B399));
  sky130_fd_sc_hd__clkbuf_4 T2Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4322));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R0_INV_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4358));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R1_INV_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R2_INV_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R2_INV_1 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4394));
  sky130_fd_sc_hd__clkbuf_4 T2Y41__R0_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4430));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R0_INV_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4466));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R1_INV_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R2_INV_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R2_INV_1 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4502));
  sky130_fd_sc_hd__clkbuf_4 T2Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4538));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R0_INV_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y42__R1_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4574));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R1_INV_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R2_INV_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R2_INV_1 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4610));
  sky130_fd_sc_hd__clkbuf_4 T2Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4646));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R0_INV_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4682));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R1_INV_0 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R2_INV_0 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R2_INV_1 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y43__R3_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4718));
  sky130_fd_sc_hd__clkbuf_4 T2Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4754));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R0_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4790));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R1_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R2_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R2_INV_1 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4826));
  sky130_fd_sc_hd__clkbuf_4 T2Y45__R0_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4862));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R0_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4898));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R1_INV_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R2_INV_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R2_INV_1 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4934));
  sky130_fd_sc_hd__clkbuf_4 T2Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4970));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R0_INV_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y46__R1_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5006));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R1_INV_0 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R2_INV_0 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R2_INV_1 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5042));
  sky130_fd_sc_hd__clkbuf_4 T2Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5078));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R0_INV_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5114));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R1_INV_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R2_INV_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R2_INV_1 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y47__R3_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5150));
  sky130_fd_sc_hd__clkbuf_4 T2Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5186));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R0_INV_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5222));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R1_INV_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R2_INV_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R2_INV_1 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5258));
  sky130_fd_sc_hd__clkbuf_4 T2Y49__R0_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5294));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R0_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5330));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R1_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R2_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R2_INV_1 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5366));
  sky130_fd_sc_hd__clkbuf_4 T2Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B435));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R0_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B471));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R1_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R2_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R2_INV_1 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B507));
  sky130_fd_sc_hd__clkbuf_4 T2Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5402));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R0_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y50__R1_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5438));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R1_INV_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R2_INV_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R2_INV_1 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5474));
  sky130_fd_sc_hd__clkbuf_4 T2Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5510));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R0_INV_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5546));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R1_INV_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R2_INV_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R2_INV_1 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y51__R3_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5582));
  sky130_fd_sc_hd__clkbuf_4 T2Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5618));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R0_INV_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5654));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R1_INV_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R2_INV_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R2_INV_1 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5690));
  sky130_fd_sc_hd__clkbuf_4 T2Y53__R0_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5726));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R0_INV_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5762));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R1_INV_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R2_INV_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R2_INV_1 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5798));
  sky130_fd_sc_hd__clkbuf_4 T2Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5834));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R0_INV_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y54__R1_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5870));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R1_INV_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R2_INV_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R2_INV_1 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5906));
  sky130_fd_sc_hd__clkbuf_4 T2Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5942));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R0_INV_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5978));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R1_INV_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R2_INV_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R2_INV_1 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y55__R3_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6014));
  sky130_fd_sc_hd__clkbuf_4 T2Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6050));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R0_INV_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6086));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R1_INV_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R2_INV_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R2_INV_1 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6122));
  sky130_fd_sc_hd__clkbuf_4 T2Y57__R0_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6158));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R0_INV_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6194));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R1_INV_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R2_INV_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R2_INV_1 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6230));
  sky130_fd_sc_hd__clkbuf_4 T2Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6266));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R0_INV_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y58__R1_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6302));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R1_INV_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R2_INV_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R2_INV_1 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6338));
  sky130_fd_sc_hd__clkbuf_4 T2Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6374));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R0_INV_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6410));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R1_INV_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R2_INV_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R2_INV_1 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y59__R3_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6446));
  sky130_fd_sc_hd__clkbuf_4 T2Y5__R0_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B543));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R0_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B579));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R1_INV_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R2_INV_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R2_INV_1 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B615));
  sky130_fd_sc_hd__clkbuf_4 T2Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6482));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R0_INV_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6518));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R1_INV_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R2_INV_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R2_INV_1 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6554));
  sky130_fd_sc_hd__clkbuf_4 T2Y61__R0_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6590));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R0_INV_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6626));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R1_INV_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R2_INV_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R2_INV_1 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6662));
  sky130_fd_sc_hd__clkbuf_4 T2Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6698));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R0_INV_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y62__R1_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6734));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R1_INV_0 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R2_INV_0 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R2_INV_1 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6770));
  sky130_fd_sc_hd__clkbuf_4 T2Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6806));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R0_INV_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6842));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R1_INV_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R2_INV_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R2_INV_1 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y63__R3_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6878));
  sky130_fd_sc_hd__clkbuf_4 T2Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6914));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R0_INV_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6950));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R1_INV_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R2_INV_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R2_INV_1 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6986));
  sky130_fd_sc_hd__clkbuf_4 T2Y65__R0_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7022));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R0_INV_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7058));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R1_INV_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R2_INV_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R2_INV_1 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7094));
  sky130_fd_sc_hd__clkbuf_4 T2Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7130));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R0_INV_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y66__R1_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7166));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R1_INV_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R2_INV_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R2_INV_1 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7202));
  sky130_fd_sc_hd__clkbuf_4 T2Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7238));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R0_INV_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7274));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R1_INV_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R2_INV_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R2_INV_1 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y67__R3_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7310));
  sky130_fd_sc_hd__clkbuf_4 T2Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7346));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R0_INV_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7382));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R1_INV_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R2_INV_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R2_INV_1 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7418));
  sky130_fd_sc_hd__clkbuf_4 T2Y69__R0_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7454));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R0_INV_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7490));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R1_INV_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R2_INV_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R2_INV_1 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7526));
  sky130_fd_sc_hd__clkbuf_4 T2Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B651));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R0_INV_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y6__R1_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B687));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R1_INV_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R2_INV_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R2_INV_1 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B723));
  sky130_fd_sc_hd__clkbuf_4 T2Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7562));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R0_INV_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y70__R1_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7598));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R1_INV_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R2_INV_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R2_INV_1 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7634));
  sky130_fd_sc_hd__clkbuf_4 T2Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7670));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R0_INV_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7706));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R1_INV_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R2_INV_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R2_INV_1 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y71__R3_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7742));
  sky130_fd_sc_hd__clkbuf_4 T2Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7778));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R0_INV_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7814));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R1_INV_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R2_INV_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R2_INV_1 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7850));
  sky130_fd_sc_hd__clkbuf_4 T2Y73__R0_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7886));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R0_INV_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7922));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R1_INV_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R2_INV_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R2_INV_1 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7958));
  sky130_fd_sc_hd__clkbuf_4 T2Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7994));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R0_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y74__R1_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8030));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R1_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R2_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R2_INV_1 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8066));
  sky130_fd_sc_hd__clkbuf_4 T2Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8102));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R0_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8138));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R1_INV_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R2_INV_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R2_INV_1 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y75__R3_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8174));
  sky130_fd_sc_hd__clkbuf_4 T2Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8210));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R0_INV_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8246));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R1_INV_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R2_INV_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R2_INV_1 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8282));
  sky130_fd_sc_hd__clkbuf_4 T2Y77__R0_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8318));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R0_INV_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8354));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R1_INV_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R2_INV_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R2_INV_1 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8390));
  sky130_fd_sc_hd__clkbuf_4 T2Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8426));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R0_INV_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y78__R1_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8462));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R1_INV_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R2_INV_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R2_INV_1 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8498));
  sky130_fd_sc_hd__clkbuf_4 T2Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8534));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R0_INV_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8570));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R1_INV_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R2_INV_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R2_INV_1 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y79__R3_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8606));
  sky130_fd_sc_hd__clkbuf_4 T2Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B759));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R0_INV_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B795));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R1_INV_0 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R2_INV_0 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R2_INV_1 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y7__R3_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B831));
  sky130_fd_sc_hd__clkbuf_4 T2Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8642));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R0_INV_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8678));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R1_INV_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R2_INV_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R2_INV_1 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8714));
  sky130_fd_sc_hd__clkbuf_4 T2Y81__R0_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8750));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R0_INV_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8786));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R1_INV_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R2_INV_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R2_INV_1 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8822));
  sky130_fd_sc_hd__clkbuf_4 T2Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8858));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R0_INV_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y82__R1_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8894));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R1_INV_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R2_INV_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R2_INV_1 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8930));
  sky130_fd_sc_hd__clkbuf_4 T2Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8966));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R0_INV_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9002));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R1_INV_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R2_INV_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R2_INV_1 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y83__R3_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9038));
  sky130_fd_sc_hd__clkbuf_4 T2Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9074));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R0_INV_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9110));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R1_INV_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R2_INV_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R2_INV_1 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9146));
  sky130_fd_sc_hd__clkbuf_4 T2Y85__R0_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9182));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R0_INV_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9218));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R1_INV_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R2_INV_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R2_INV_1 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9254));
  sky130_fd_sc_hd__clkbuf_4 T2Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9290));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R0_INV_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y86__R1_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9326));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R1_INV_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R2_INV_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R2_INV_1 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9362));
  sky130_fd_sc_hd__clkbuf_4 T2Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9398));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R0_INV_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9434));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R1_INV_0 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R2_INV_0 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R2_INV_1 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y87__R3_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9470));
  sky130_fd_sc_hd__clkbuf_4 T2Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9506));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R0_INV_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9542));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R1_INV_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R2_INV_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R2_INV_1 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9578));
  sky130_fd_sc_hd__clkbuf_4 T2Y89__R0_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9614));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R0_INV_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9650));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R1_INV_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R2_INV_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R2_INV_1 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9686));
  sky130_fd_sc_hd__clkbuf_4 T2Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B867));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R0_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B903));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R1_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R2_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R2_INV_1 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B939));
  sky130_fd_sc_hd__clkbuf_4 T2Y9__R0_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B975));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R0_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1011));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R1_INV_0 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R2_INV_0 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R2_INV_1 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1047));
  sky130_fd_sc_hd__clkbuf_4 T30Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B40));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R0_INV_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B75));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R1_INV_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R2_INV_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R2_INV_1 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B110));
  sky130_fd_sc_hd__clkbuf_4 T30Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1111));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R0_INV_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1147));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R1_INV_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R2_INV_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R2_INV_1 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y10__R3_BUF_0 (.A(clk_L1_B73), .X(clk_L0_B1183));
  sky130_fd_sc_hd__clkbuf_4 T30Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1219));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R0_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1255));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R1_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R2_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R2_INV_1 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1291));
  sky130_fd_sc_hd__clkbuf_4 T30Y12__R0_BUF_0 (.A(clk_L1_B82), .X(clk_L0_B1327));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R0_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1363));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R1_INV_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R2_INV_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R2_INV_1 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1399));
  sky130_fd_sc_hd__clkbuf_4 T30Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1435));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R0_INV_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y13__R1_BUF_0 (.A(clk_L1_B91), .X(clk_L0_B1471));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R1_INV_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R2_INV_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R2_INV_1 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1507));
  sky130_fd_sc_hd__clkbuf_4 T30Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1543));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R0_INV_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1578));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R1_INV_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R2_INV_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R2_INV_1 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1614));
  sky130_fd_sc_hd__clkbuf_4 T30Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1650));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R0_INV_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1686));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R1_INV_0 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R2_INV_0 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R2_INV_1 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1722));
  sky130_fd_sc_hd__clkbuf_4 T30Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1758));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R0_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1794));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R1_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R2_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R2_INV_1 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1830));
  sky130_fd_sc_hd__clkbuf_4 T30Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1866));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R0_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1902));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R1_INV_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R2_INV_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R2_INV_1 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1938));
  sky130_fd_sc_hd__clkbuf_4 T30Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1974));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R0_INV_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2010));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R1_INV_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R2_INV_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R2_INV_1 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2046));
  sky130_fd_sc_hd__clkbuf_4 T30Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2082));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R0_INV_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2118));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R1_INV_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R2_INV_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R2_INV_1 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2154));
  sky130_fd_sc_hd__clkbuf_4 T30Y1__R0_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B145));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R0_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B180));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R1_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R2_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R2_INV_1 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B215));
  sky130_fd_sc_hd__clkbuf_4 T30Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2190));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R0_INV_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2226));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R1_INV_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R2_INV_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R2_INV_1 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2262));
  sky130_fd_sc_hd__clkbuf_4 T30Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2298));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R0_INV_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2334));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R1_INV_0 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R2_INV_0 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R2_INV_1 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2370));
  sky130_fd_sc_hd__clkbuf_4 T30Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2406));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R0_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2442));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R1_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R2_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R2_INV_1 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2478));
  sky130_fd_sc_hd__clkbuf_4 T30Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2514));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R0_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2550));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R1_INV_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R2_INV_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R2_INV_1 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2586));
  sky130_fd_sc_hd__clkbuf_4 T30Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2622));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R0_INV_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2658));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R1_INV_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R2_INV_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R2_INV_1 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2694));
  sky130_fd_sc_hd__clkbuf_4 T30Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2730));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R0_INV_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2766));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R1_INV_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R2_INV_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R2_INV_1 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2802));
  sky130_fd_sc_hd__clkbuf_4 T30Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2838));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R0_INV_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2874));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R1_INV_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R2_INV_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R2_INV_1 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2910));
  sky130_fd_sc_hd__clkbuf_4 T30Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2946));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R0_INV_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2982));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R1_INV_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R2_INV_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R2_INV_1 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3018));
  sky130_fd_sc_hd__clkbuf_4 T30Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3054));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R0_INV_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3090));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R1_INV_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R2_INV_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R2_INV_1 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3126));
  sky130_fd_sc_hd__clkbuf_4 T30Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3162));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R0_INV_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3198));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R1_INV_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R2_INV_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R2_INV_1 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3234));
  sky130_fd_sc_hd__clkbuf_4 T30Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B250));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R0_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B285));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R1_INV_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R2_INV_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R2_INV_1 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y2__R3_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B321));
  sky130_fd_sc_hd__clkbuf_4 T30Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3270));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R0_INV_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3306));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R1_INV_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R2_INV_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R2_INV_1 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3342));
  sky130_fd_sc_hd__clkbuf_4 T30Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3378));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R0_INV_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3414));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R1_INV_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R2_INV_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R2_INV_1 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3450));
  sky130_fd_sc_hd__clkbuf_4 T30Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3486));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R0_INV_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3522));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R1_INV_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R2_INV_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R2_INV_1 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3558));
  sky130_fd_sc_hd__clkbuf_4 T30Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3594));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R0_INV_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3630));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R1_INV_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R2_INV_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R2_INV_1 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3666));
  sky130_fd_sc_hd__clkbuf_4 T30Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3702));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R0_INV_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3738));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R1_INV_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R2_INV_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R2_INV_1 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3774));
  sky130_fd_sc_hd__clkbuf_4 T30Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3810));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R0_INV_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3846));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R1_INV_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R2_INV_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R2_INV_1 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3882));
  sky130_fd_sc_hd__clkbuf_4 T30Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3918));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R0_INV_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3954));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R1_INV_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R2_INV_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R2_INV_1 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3990));
  sky130_fd_sc_hd__clkbuf_4 T30Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4026));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R0_INV_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4062));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R1_INV_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R2_INV_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R2_INV_1 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4098));
  sky130_fd_sc_hd__clkbuf_4 T30Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4134));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R0_INV_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4170));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R1_INV_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R2_INV_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R2_INV_1 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4206));
  sky130_fd_sc_hd__clkbuf_4 T30Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4242));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R0_INV_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4278));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R1_INV_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R2_INV_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R2_INV_1 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4314));
  sky130_fd_sc_hd__clkbuf_4 T30Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B356));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R0_INV_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B391));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R1_INV_0 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R2_INV_0 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R2_INV_1 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B427));
  sky130_fd_sc_hd__clkbuf_4 T30Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4350));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R0_INV_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4386));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R1_INV_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R2_INV_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R2_INV_1 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4422));
  sky130_fd_sc_hd__clkbuf_4 T30Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4458));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R0_INV_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4494));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R1_INV_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R2_INV_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R2_INV_1 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4530));
  sky130_fd_sc_hd__clkbuf_4 T30Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4566));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R0_INV_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4602));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R1_INV_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R2_INV_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R2_INV_1 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4638));
  sky130_fd_sc_hd__clkbuf_4 T30Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4674));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R0_INV_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4710));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R1_INV_0 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R2_INV_0 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R2_INV_1 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4746));
  sky130_fd_sc_hd__clkbuf_4 T30Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4782));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R0_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4818));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R1_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R2_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R2_INV_1 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4854));
  sky130_fd_sc_hd__clkbuf_4 T30Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4890));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R0_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4926));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R1_INV_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R2_INV_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R2_INV_1 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4962));
  sky130_fd_sc_hd__clkbuf_4 T30Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4998));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R0_INV_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5034));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R1_INV_0 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R2_INV_0 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R2_INV_1 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5070));
  sky130_fd_sc_hd__clkbuf_4 T30Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5106));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R0_INV_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5142));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R1_INV_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R2_INV_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R2_INV_1 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5178));
  sky130_fd_sc_hd__clkbuf_4 T30Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5214));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R0_INV_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5250));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R1_INV_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R2_INV_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R2_INV_1 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5286));
  sky130_fd_sc_hd__clkbuf_4 T30Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5322));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R0_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5358));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R1_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R2_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R2_INV_1 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5394));
  sky130_fd_sc_hd__clkbuf_4 T30Y4__R0_BUF_0 (.A(clk_L1_B28), .X(clk_L0_B463));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R0_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B499));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R1_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R2_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R2_INV_1 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B535));
  sky130_fd_sc_hd__clkbuf_4 T30Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5430));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R0_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5466));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R1_INV_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R2_INV_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R2_INV_1 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5502));
  sky130_fd_sc_hd__clkbuf_4 T30Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5538));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R0_INV_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5574));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R1_INV_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R2_INV_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R2_INV_1 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5610));
  sky130_fd_sc_hd__clkbuf_4 T30Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5646));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R0_INV_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5682));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R1_INV_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R2_INV_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R2_INV_1 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5718));
  sky130_fd_sc_hd__clkbuf_4 T30Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5754));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R0_INV_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5790));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R1_INV_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R2_INV_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R2_INV_1 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5826));
  sky130_fd_sc_hd__clkbuf_4 T30Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5862));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R0_INV_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5898));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R1_INV_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R2_INV_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R2_INV_1 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5934));
  sky130_fd_sc_hd__clkbuf_4 T30Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5970));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R0_INV_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6006));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R1_INV_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R2_INV_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R2_INV_1 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6042));
  sky130_fd_sc_hd__clkbuf_4 T30Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6078));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R0_INV_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6114));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R1_INV_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R2_INV_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R2_INV_1 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6150));
  sky130_fd_sc_hd__clkbuf_4 T30Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6186));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R0_INV_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6222));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R1_INV_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R2_INV_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R2_INV_1 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6258));
  sky130_fd_sc_hd__clkbuf_4 T30Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6294));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R0_INV_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6330));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R1_INV_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R2_INV_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R2_INV_1 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6366));
  sky130_fd_sc_hd__clkbuf_4 T30Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6402));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R0_INV_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6438));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R1_INV_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R2_INV_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R2_INV_1 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6474));
  sky130_fd_sc_hd__clkbuf_4 T30Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B571));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R0_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y5__R1_BUF_0 (.A(clk_L1_B37), .X(clk_L0_B607));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R1_INV_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R2_INV_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R2_INV_1 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B643));
  sky130_fd_sc_hd__clkbuf_4 T30Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6510));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R0_INV_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6546));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R1_INV_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R2_INV_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R2_INV_1 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6582));
  sky130_fd_sc_hd__clkbuf_4 T30Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6618));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R0_INV_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6654));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R1_INV_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R2_INV_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R2_INV_1 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6690));
  sky130_fd_sc_hd__clkbuf_4 T30Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6726));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R0_INV_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6762));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R1_INV_0 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R2_INV_0 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R2_INV_1 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6798));
  sky130_fd_sc_hd__clkbuf_4 T30Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6834));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R0_INV_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6870));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R1_INV_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R2_INV_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R2_INV_1 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6906));
  sky130_fd_sc_hd__clkbuf_4 T30Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6942));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R0_INV_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6978));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R1_INV_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R2_INV_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R2_INV_1 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7014));
  sky130_fd_sc_hd__clkbuf_4 T30Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7050));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R0_INV_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7086));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R1_INV_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R2_INV_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R2_INV_1 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7122));
  sky130_fd_sc_hd__clkbuf_4 T30Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7158));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R0_INV_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7194));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R1_INV_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R2_INV_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R2_INV_1 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7230));
  sky130_fd_sc_hd__clkbuf_4 T30Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7266));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R0_INV_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7302));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R1_INV_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R2_INV_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R2_INV_1 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7338));
  sky130_fd_sc_hd__clkbuf_4 T30Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7374));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R0_INV_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7410));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R1_INV_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R2_INV_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R2_INV_1 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7446));
  sky130_fd_sc_hd__clkbuf_4 T30Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7482));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R0_INV_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7518));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R1_INV_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R2_INV_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R2_INV_1 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7554));
  sky130_fd_sc_hd__clkbuf_4 T30Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B679));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R0_INV_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B715));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R1_INV_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R2_INV_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R2_INV_1 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y6__R3_BUF_0 (.A(clk_L1_B46), .X(clk_L0_B751));
  sky130_fd_sc_hd__clkbuf_4 T30Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7590));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R0_INV_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7626));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R1_INV_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R2_INV_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R2_INV_1 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7662));
  sky130_fd_sc_hd__clkbuf_4 T30Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7698));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R0_INV_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7734));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R1_INV_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R2_INV_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R2_INV_1 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7770));
  sky130_fd_sc_hd__clkbuf_4 T30Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7806));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R0_INV_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7842));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R1_INV_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R2_INV_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R2_INV_1 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7878));
  sky130_fd_sc_hd__clkbuf_4 T30Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7914));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R0_INV_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7950));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R1_INV_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R2_INV_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R2_INV_1 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7986));
  sky130_fd_sc_hd__clkbuf_4 T30Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8022));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R0_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8058));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R1_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R2_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R2_INV_1 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8094));
  sky130_fd_sc_hd__clkbuf_4 T30Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8130));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R0_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8166));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R1_INV_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R2_INV_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R2_INV_1 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8202));
  sky130_fd_sc_hd__clkbuf_4 T30Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8238));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R0_INV_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8274));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R1_INV_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R2_INV_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R2_INV_1 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8310));
  sky130_fd_sc_hd__clkbuf_4 T30Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8346));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R0_INV_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8382));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R1_INV_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R2_INV_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R2_INV_1 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8418));
  sky130_fd_sc_hd__clkbuf_4 T30Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8454));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R0_INV_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8490));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R1_INV_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R2_INV_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R2_INV_1 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8526));
  sky130_fd_sc_hd__clkbuf_4 T30Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8562));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R0_INV_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8598));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R1_INV_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R2_INV_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R2_INV_1 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8634));
  sky130_fd_sc_hd__clkbuf_4 T30Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B787));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R0_INV_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B823));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R1_INV_0 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R2_INV_0 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R2_INV_1 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B859));
  sky130_fd_sc_hd__clkbuf_4 T30Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8670));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R0_INV_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8706));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R1_INV_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R2_INV_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R2_INV_1 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8742));
  sky130_fd_sc_hd__clkbuf_4 T30Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8778));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R0_INV_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8814));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R1_INV_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R2_INV_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R2_INV_1 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8850));
  sky130_fd_sc_hd__clkbuf_4 T30Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8886));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R0_INV_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8922));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R1_INV_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R2_INV_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R2_INV_1 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8958));
  sky130_fd_sc_hd__clkbuf_4 T30Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8994));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R0_INV_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9030));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R1_INV_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R2_INV_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R2_INV_1 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9066));
  sky130_fd_sc_hd__clkbuf_4 T30Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9102));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R0_INV_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9138));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R1_INV_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R2_INV_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R2_INV_1 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9174));
  sky130_fd_sc_hd__clkbuf_4 T30Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9210));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R0_INV_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9246));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R1_INV_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R2_INV_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R2_INV_1 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9282));
  sky130_fd_sc_hd__clkbuf_4 T30Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9318));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R0_INV_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9354));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R1_INV_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R2_INV_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R2_INV_1 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9390));
  sky130_fd_sc_hd__clkbuf_4 T30Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9426));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R0_INV_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9462));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R1_INV_0 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R2_INV_0 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R2_INV_1 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9498));
  sky130_fd_sc_hd__clkbuf_4 T30Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9534));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R0_INV_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9570));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R1_INV_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R2_INV_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R2_INV_1 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9606));
  sky130_fd_sc_hd__clkbuf_4 T30Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9642));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R0_INV_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9678));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R1_INV_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R2_INV_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R2_INV_1 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9714));
  sky130_fd_sc_hd__clkbuf_4 T30Y8__R0_BUF_0 (.A(clk_L1_B55), .X(clk_L0_B895));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R0_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B931));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R1_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R2_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R2_INV_1 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B967));
  sky130_fd_sc_hd__clkbuf_4 T30Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1003));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R0_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y9__R1_BUF_0 (.A(clk_L1_B64), .X(clk_L0_B1039));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R1_INV_0 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R2_INV_0 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R2_INV_1 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1075));
  sky130_fd_sc_hd__clkbuf_4 T31Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B41));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R0_INV_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B76));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R1_INV_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R2_INV_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R2_INV_1 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y0__R3_BUF_0 (.A(clk_L1_B6), .X(clk_L0_B111));
  sky130_fd_sc_hd__clkbuf_4 T31Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1112));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R0_INV_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1148));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R1_INV_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R2_INV_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R2_INV_1 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y10__R3_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B74));
  sky130_fd_sc_hd__clkbuf_4 T31Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1220));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R0_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1256));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R1_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R2_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R2_INV_1 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1292));
  sky130_fd_sc_hd__clkbuf_4 T31Y12__R0_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B83));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R0_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1364));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R1_INV_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R2_INV_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R2_INV_1 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1400));
  sky130_fd_sc_hd__clkbuf_4 T31Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1436));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R0_INV_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y13__R1_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B92));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R1_INV_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R2_INV_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R2_INV_1 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1508));
  sky130_fd_sc_hd__clkbuf_4 T31Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1544));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R0_INV_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1579));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R1_INV_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R2_INV_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R2_INV_1 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y14__R3_BUF_0 (.A(clk_L1_B100), .X(clk_L0_B1615));
  sky130_fd_sc_hd__clkbuf_4 T31Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1651));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R0_INV_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1687));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R1_INV_0 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R2_INV_0 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R2_INV_1 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1723));
  sky130_fd_sc_hd__clkbuf_4 T31Y16__R0_BUF_0 (.A(clk_L1_B109), .X(clk_L0_B1759));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R0_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1795));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R1_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R2_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R2_INV_1 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1831));
  sky130_fd_sc_hd__clkbuf_4 T31Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1867));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R0_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y17__R1_BUF_0 (.A(clk_L1_B118), .X(clk_L0_B1903));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R1_INV_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R2_INV_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R2_INV_1 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1939));
  sky130_fd_sc_hd__clkbuf_4 T31Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1975));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R0_INV_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2011));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R1_INV_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R2_INV_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R2_INV_1 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y18__R3_BUF_0 (.A(clk_L1_B127), .X(clk_L0_B2047));
  sky130_fd_sc_hd__clkbuf_4 T31Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2083));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R0_INV_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2119));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R1_INV_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R2_INV_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R2_INV_1 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2155));
  sky130_fd_sc_hd__clkbuf_4 T31Y1__R0_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B146));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R0_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B181));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R1_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R2_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R2_INV_1 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B216));
  sky130_fd_sc_hd__clkbuf_4 T31Y20__R0_BUF_0 (.A(clk_L1_B136), .X(clk_L0_B2191));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R0_INV_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2227));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R1_INV_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R2_INV_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R2_INV_1 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2263));
  sky130_fd_sc_hd__clkbuf_4 T31Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2299));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R0_INV_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y21__R1_BUF_0 (.A(clk_L1_B145), .X(clk_L0_B2335));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R1_INV_0 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R2_INV_0 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R2_INV_1 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2371));
  sky130_fd_sc_hd__clkbuf_4 T31Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2407));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R0_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2443));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R1_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R2_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R2_INV_1 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y22__R3_BUF_0 (.A(clk_L1_B154), .X(clk_L0_B2479));
  sky130_fd_sc_hd__clkbuf_4 T31Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2515));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R0_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2551));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R1_INV_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R2_INV_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R2_INV_1 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2587));
  sky130_fd_sc_hd__clkbuf_4 T31Y24__R0_BUF_0 (.A(clk_L1_B163), .X(clk_L0_B2623));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R0_INV_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2659));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R1_INV_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R2_INV_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R2_INV_1 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2695));
  sky130_fd_sc_hd__clkbuf_4 T31Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2731));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R0_INV_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y25__R1_BUF_0 (.A(clk_L1_B172), .X(clk_L0_B2767));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R1_INV_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R2_INV_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R2_INV_1 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2803));
  sky130_fd_sc_hd__clkbuf_4 T31Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2839));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R0_INV_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2875));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R1_INV_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R2_INV_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R2_INV_1 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y26__R3_BUF_0 (.A(clk_L1_B181), .X(clk_L0_B2911));
  sky130_fd_sc_hd__clkbuf_4 T31Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2947));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R0_INV_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2983));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R1_INV_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R2_INV_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R2_INV_1 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3019));
  sky130_fd_sc_hd__clkbuf_4 T31Y28__R0_BUF_0 (.A(clk_L1_B190), .X(clk_L0_B3055));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R0_INV_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3091));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R1_INV_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R2_INV_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R2_INV_1 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3127));
  sky130_fd_sc_hd__clkbuf_4 T31Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3163));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R0_INV_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y29__R1_BUF_0 (.A(clk_L1_B199), .X(clk_L0_B3199));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R1_INV_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R2_INV_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R2_INV_1 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3235));
  sky130_fd_sc_hd__clkbuf_4 T31Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B251));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R0_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B286));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R1_INV_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R2_INV_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R2_INV_1 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y2__R3_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B322));
  sky130_fd_sc_hd__clkbuf_4 T31Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3271));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R0_INV_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3307));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R1_INV_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R2_INV_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R2_INV_1 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y30__R3_BUF_0 (.A(clk_L1_B208), .X(clk_L0_B3343));
  sky130_fd_sc_hd__clkbuf_4 T31Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3379));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R0_INV_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3415));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R1_INV_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R2_INV_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R2_INV_1 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3451));
  sky130_fd_sc_hd__clkbuf_4 T31Y32__R0_BUF_0 (.A(clk_L1_B217), .X(clk_L0_B3487));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R0_INV_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3523));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R1_INV_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R2_INV_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R2_INV_1 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3559));
  sky130_fd_sc_hd__clkbuf_4 T31Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3595));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R0_INV_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y33__R1_BUF_0 (.A(clk_L1_B226), .X(clk_L0_B3631));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R1_INV_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R2_INV_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R2_INV_1 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3667));
  sky130_fd_sc_hd__clkbuf_4 T31Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3703));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R0_INV_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3739));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R1_INV_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R2_INV_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R2_INV_1 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y34__R3_BUF_0 (.A(clk_L1_B235), .X(clk_L0_B3775));
  sky130_fd_sc_hd__clkbuf_4 T31Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3811));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R0_INV_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3847));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R1_INV_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R2_INV_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R2_INV_1 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3883));
  sky130_fd_sc_hd__clkbuf_4 T31Y36__R0_BUF_0 (.A(clk_L1_B244), .X(clk_L0_B3919));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R0_INV_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3955));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R1_INV_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R2_INV_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R2_INV_1 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3991));
  sky130_fd_sc_hd__clkbuf_4 T31Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4027));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R0_INV_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y37__R1_BUF_0 (.A(clk_L1_B253), .X(clk_L0_B4063));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R1_INV_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R2_INV_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R2_INV_1 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4099));
  sky130_fd_sc_hd__clkbuf_4 T31Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4135));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R0_INV_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4171));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R1_INV_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R2_INV_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R2_INV_1 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y38__R3_BUF_0 (.A(clk_L1_B262), .X(clk_L0_B4207));
  sky130_fd_sc_hd__clkbuf_4 T31Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4243));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R0_INV_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4279));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R1_INV_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R2_INV_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R2_INV_1 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4315));
  sky130_fd_sc_hd__clkbuf_4 T31Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B357));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R0_INV_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B392));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R1_INV_0 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R2_INV_0 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R2_INV_1 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B428));
  sky130_fd_sc_hd__clkbuf_4 T31Y40__R0_BUF_0 (.A(clk_L1_B271), .X(clk_L0_B4351));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R0_INV_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4387));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R1_INV_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R2_INV_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R2_INV_1 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4423));
  sky130_fd_sc_hd__clkbuf_4 T31Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4459));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R0_INV_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y41__R1_BUF_0 (.A(clk_L1_B280), .X(clk_L0_B4495));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R1_INV_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R2_INV_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R2_INV_1 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4531));
  sky130_fd_sc_hd__clkbuf_4 T31Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4567));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R0_INV_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4603));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R1_INV_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R2_INV_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R2_INV_1 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y42__R3_BUF_0 (.A(clk_L1_B289), .X(clk_L0_B4639));
  sky130_fd_sc_hd__clkbuf_4 T31Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4675));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R0_INV_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4711));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R1_INV_0 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R2_INV_0 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R2_INV_1 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4747));
  sky130_fd_sc_hd__clkbuf_4 T31Y44__R0_BUF_0 (.A(clk_L1_B298), .X(clk_L0_B4783));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R0_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4819));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R1_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R2_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R2_INV_1 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4855));
  sky130_fd_sc_hd__clkbuf_4 T31Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4891));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R0_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y45__R1_BUF_0 (.A(clk_L1_B307), .X(clk_L0_B4927));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R1_INV_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R2_INV_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R2_INV_1 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4963));
  sky130_fd_sc_hd__clkbuf_4 T31Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B4999));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R0_INV_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5035));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R1_INV_0 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R2_INV_0 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R2_INV_1 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y46__R3_BUF_0 (.A(clk_L1_B316), .X(clk_L0_B5071));
  sky130_fd_sc_hd__clkbuf_4 T31Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5107));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R0_INV_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5143));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R1_INV_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R2_INV_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R2_INV_1 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5179));
  sky130_fd_sc_hd__clkbuf_4 T31Y48__R0_BUF_0 (.A(clk_L1_B325), .X(clk_L0_B5215));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R0_INV_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5251));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R1_INV_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R2_INV_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R2_INV_1 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5287));
  sky130_fd_sc_hd__clkbuf_4 T31Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5323));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R0_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y49__R1_BUF_0 (.A(clk_L1_B334), .X(clk_L0_B5359));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R1_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R2_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R2_INV_1 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5395));
  sky130_fd_sc_hd__clkbuf_4 T31Y4__R0_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B29));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R0_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B500));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R1_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R2_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R2_INV_1 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B536));
  sky130_fd_sc_hd__clkbuf_4 T31Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5431));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R0_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5467));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R1_INV_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R2_INV_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R2_INV_1 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y50__R3_BUF_0 (.A(clk_L1_B343), .X(clk_L0_B5503));
  sky130_fd_sc_hd__clkbuf_4 T31Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5539));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R0_INV_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5575));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R1_INV_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R2_INV_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R2_INV_1 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5611));
  sky130_fd_sc_hd__clkbuf_4 T31Y52__R0_BUF_0 (.A(clk_L1_B352), .X(clk_L0_B5647));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R0_INV_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5683));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R1_INV_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R2_INV_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R2_INV_1 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5719));
  sky130_fd_sc_hd__clkbuf_4 T31Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5755));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R0_INV_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y53__R1_BUF_0 (.A(clk_L1_B361), .X(clk_L0_B5791));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R1_INV_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R2_INV_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R2_INV_1 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5827));
  sky130_fd_sc_hd__clkbuf_4 T31Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5863));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R0_INV_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5899));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R1_INV_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R2_INV_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R2_INV_1 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y54__R3_BUF_0 (.A(clk_L1_B370), .X(clk_L0_B5935));
  sky130_fd_sc_hd__clkbuf_4 T31Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5971));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R0_INV_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6007));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R1_INV_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R2_INV_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R2_INV_1 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6043));
  sky130_fd_sc_hd__clkbuf_4 T31Y56__R0_BUF_0 (.A(clk_L1_B379), .X(clk_L0_B6079));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R0_INV_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6115));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R1_INV_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R2_INV_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R2_INV_1 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6151));
  sky130_fd_sc_hd__clkbuf_4 T31Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6187));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R0_INV_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y57__R1_BUF_0 (.A(clk_L1_B388), .X(clk_L0_B6223));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R1_INV_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R2_INV_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R2_INV_1 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6259));
  sky130_fd_sc_hd__clkbuf_4 T31Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6295));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R0_INV_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6331));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R1_INV_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R2_INV_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R2_INV_1 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y58__R3_BUF_0 (.A(clk_L1_B397), .X(clk_L0_B6367));
  sky130_fd_sc_hd__clkbuf_4 T31Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6403));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R0_INV_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6439));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R1_INV_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R2_INV_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R2_INV_1 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6475));
  sky130_fd_sc_hd__clkbuf_4 T31Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B572));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R0_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y5__R1_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B38));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R1_INV_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R2_INV_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R2_INV_1 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B644));
  sky130_fd_sc_hd__clkbuf_4 T31Y60__R0_BUF_0 (.A(clk_L1_B406), .X(clk_L0_B6511));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R0_INV_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6547));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R1_INV_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R2_INV_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R2_INV_1 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6583));
  sky130_fd_sc_hd__clkbuf_4 T31Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6619));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R0_INV_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y61__R1_BUF_0 (.A(clk_L1_B415), .X(clk_L0_B6655));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R1_INV_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R2_INV_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R2_INV_1 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6691));
  sky130_fd_sc_hd__clkbuf_4 T31Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6727));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R0_INV_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6763));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R1_INV_0 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R2_INV_0 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R2_INV_1 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y62__R3_BUF_0 (.A(clk_L1_B424), .X(clk_L0_B6799));
  sky130_fd_sc_hd__clkbuf_4 T31Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6835));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R0_INV_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6871));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R1_INV_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R2_INV_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R2_INV_1 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6907));
  sky130_fd_sc_hd__clkbuf_4 T31Y64__R0_BUF_0 (.A(clk_L1_B433), .X(clk_L0_B6943));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R0_INV_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6979));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R1_INV_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R2_INV_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R2_INV_1 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7015));
  sky130_fd_sc_hd__clkbuf_4 T31Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7051));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R0_INV_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y65__R1_BUF_0 (.A(clk_L1_B442), .X(clk_L0_B7087));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R1_INV_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R2_INV_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R2_INV_1 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7123));
  sky130_fd_sc_hd__clkbuf_4 T31Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7159));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R0_INV_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7195));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R1_INV_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R2_INV_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R2_INV_1 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y66__R3_BUF_0 (.A(clk_L1_B451), .X(clk_L0_B7231));
  sky130_fd_sc_hd__clkbuf_4 T31Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7267));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R0_INV_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7303));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R1_INV_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R2_INV_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R2_INV_1 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7339));
  sky130_fd_sc_hd__clkbuf_4 T31Y68__R0_BUF_0 (.A(clk_L1_B460), .X(clk_L0_B7375));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R0_INV_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7411));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R1_INV_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R2_INV_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R2_INV_1 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7447));
  sky130_fd_sc_hd__clkbuf_4 T31Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7483));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R0_INV_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y69__R1_BUF_0 (.A(clk_L1_B469), .X(clk_L0_B7519));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R1_INV_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R2_INV_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R2_INV_1 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7555));
  sky130_fd_sc_hd__clkbuf_4 T31Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B680));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R0_INV_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B716));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R1_INV_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R2_INV_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R2_INV_1 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y6__R3_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B47));
  sky130_fd_sc_hd__clkbuf_4 T31Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7591));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R0_INV_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7627));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R1_INV_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R2_INV_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R2_INV_1 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y70__R3_BUF_0 (.A(clk_L1_B478), .X(clk_L0_B7663));
  sky130_fd_sc_hd__clkbuf_4 T31Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7699));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R0_INV_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7735));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R1_INV_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R2_INV_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R2_INV_1 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7771));
  sky130_fd_sc_hd__clkbuf_4 T31Y72__R0_BUF_0 (.A(clk_L1_B487), .X(clk_L0_B7807));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R0_INV_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7843));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R1_INV_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R2_INV_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R2_INV_1 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7879));
  sky130_fd_sc_hd__clkbuf_4 T31Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7915));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R0_INV_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y73__R1_BUF_0 (.A(clk_L1_B496), .X(clk_L0_B7951));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R1_INV_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R2_INV_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R2_INV_1 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7987));
  sky130_fd_sc_hd__clkbuf_4 T31Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8023));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R0_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8059));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R1_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R2_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R2_INV_1 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y74__R3_BUF_0 (.A(clk_L1_B505), .X(clk_L0_B8095));
  sky130_fd_sc_hd__clkbuf_4 T31Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8131));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R0_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8167));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R1_INV_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R2_INV_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R2_INV_1 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8203));
  sky130_fd_sc_hd__clkbuf_4 T31Y76__R0_BUF_0 (.A(clk_L1_B514), .X(clk_L0_B8239));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R0_INV_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8275));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R1_INV_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R2_INV_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R2_INV_1 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8311));
  sky130_fd_sc_hd__clkbuf_4 T31Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8347));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R0_INV_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y77__R1_BUF_0 (.A(clk_L1_B523), .X(clk_L0_B8383));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R1_INV_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R2_INV_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R2_INV_1 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8419));
  sky130_fd_sc_hd__clkbuf_4 T31Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8455));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R0_INV_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8491));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R1_INV_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R2_INV_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R2_INV_1 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y78__R3_BUF_0 (.A(clk_L1_B532), .X(clk_L0_B8527));
  sky130_fd_sc_hd__clkbuf_4 T31Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8563));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R0_INV_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8599));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R1_INV_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R2_INV_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R2_INV_1 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8635));
  sky130_fd_sc_hd__clkbuf_4 T31Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B788));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R0_INV_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B824));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R1_INV_0 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R2_INV_0 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R2_INV_1 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B860));
  sky130_fd_sc_hd__clkbuf_4 T31Y80__R0_BUF_0 (.A(clk_L1_B541), .X(clk_L0_B8671));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R0_INV_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8707));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R1_INV_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R2_INV_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R2_INV_1 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8743));
  sky130_fd_sc_hd__clkbuf_4 T31Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8779));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R0_INV_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y81__R1_BUF_0 (.A(clk_L1_B550), .X(clk_L0_B8815));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R1_INV_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R2_INV_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R2_INV_1 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8851));
  sky130_fd_sc_hd__clkbuf_4 T31Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8887));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R0_INV_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8923));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R1_INV_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R2_INV_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R2_INV_1 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y82__R3_BUF_0 (.A(clk_L1_B559), .X(clk_L0_B8959));
  sky130_fd_sc_hd__clkbuf_4 T31Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8995));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R0_INV_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9031));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R1_INV_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R2_INV_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R2_INV_1 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9067));
  sky130_fd_sc_hd__clkbuf_4 T31Y84__R0_BUF_0 (.A(clk_L1_B568), .X(clk_L0_B9103));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R0_INV_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9139));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R1_INV_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R2_INV_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R2_INV_1 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9175));
  sky130_fd_sc_hd__clkbuf_4 T31Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9211));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R0_INV_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y85__R1_BUF_0 (.A(clk_L1_B577), .X(clk_L0_B9247));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R1_INV_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R2_INV_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R2_INV_1 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9283));
  sky130_fd_sc_hd__clkbuf_4 T31Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9319));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R0_INV_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9355));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R1_INV_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R2_INV_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R2_INV_1 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y86__R3_BUF_0 (.A(clk_L1_B586), .X(clk_L0_B9391));
  sky130_fd_sc_hd__clkbuf_4 T31Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9427));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R0_INV_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9463));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R1_INV_0 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R2_INV_0 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R2_INV_1 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9499));
  sky130_fd_sc_hd__clkbuf_4 T31Y88__R0_BUF_0 (.A(clk_L1_B595), .X(clk_L0_B9535));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R0_INV_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9571));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R1_INV_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R2_INV_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R2_INV_1 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9607));
  sky130_fd_sc_hd__clkbuf_4 T31Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9643));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R0_INV_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y89__R1_BUF_0 (.A(clk_L1_B604), .X(clk_L0_B9679));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R1_INV_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R2_INV_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R2_INV_1 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9715));
  sky130_fd_sc_hd__clkbuf_4 T31Y8__R0_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B56));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R0_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B932));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R1_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R2_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R2_INV_1 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B968));
  sky130_fd_sc_hd__clkbuf_4 T31Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1004));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R0_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y9__R1_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B65));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R1_INV_0 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R2_INV_0 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R2_INV_1 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1076));
  sky130_fd_sc_hd__clkbuf_4 T32Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B42));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R0_INV_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B77));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R1_INV_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R2_INV_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R2_INV_1 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y0__R3_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B7));
  sky130_fd_sc_hd__clkbuf_4 T32Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1113));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R0_INV_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1149));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R1_INV_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R2_INV_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R2_INV_1 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y10__R3_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1185));
  sky130_fd_sc_hd__clkbuf_4 T32Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1221));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R0_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1257));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R1_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R2_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R2_INV_1 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1293));
  sky130_fd_sc_hd__clkbuf_4 T32Y12__R0_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1329));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R0_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1365));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R1_INV_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R2_INV_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R2_INV_1 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1401));
  sky130_fd_sc_hd__clkbuf_4 T32Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1437));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R0_INV_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y13__R1_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1473));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R1_INV_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R2_INV_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R2_INV_1 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1509));
  sky130_fd_sc_hd__clkbuf_4 T32Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1545));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R0_INV_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1580));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R1_INV_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R2_INV_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R2_INV_1 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y14__R3_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B101));
  sky130_fd_sc_hd__clkbuf_4 T32Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1652));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R0_INV_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1688));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R1_INV_0 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R2_INV_0 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R2_INV_1 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1724));
  sky130_fd_sc_hd__clkbuf_4 T32Y16__R0_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B110));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R0_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1796));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R1_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R2_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R2_INV_1 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1832));
  sky130_fd_sc_hd__clkbuf_4 T32Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1868));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R0_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y17__R1_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B119));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R1_INV_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R2_INV_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R2_INV_1 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1940));
  sky130_fd_sc_hd__clkbuf_4 T32Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1976));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R0_INV_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2012));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R1_INV_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R2_INV_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R2_INV_1 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y18__R3_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B8));
  sky130_fd_sc_hd__clkbuf_4 T32Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2084));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R0_INV_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2120));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R1_INV_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R2_INV_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R2_INV_1 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2156));
  sky130_fd_sc_hd__clkbuf_4 T32Y1__R0_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B147));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R0_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B182));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R1_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R2_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R2_INV_1 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B217));
  sky130_fd_sc_hd__clkbuf_4 T32Y20__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B137));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R0_INV_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2228));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R1_INV_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R2_INV_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R2_INV_1 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2264));
  sky130_fd_sc_hd__clkbuf_4 T32Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2300));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R0_INV_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y21__R1_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B146));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R1_INV_0 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R2_INV_0 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R2_INV_1 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2372));
  sky130_fd_sc_hd__clkbuf_4 T32Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2408));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R0_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2444));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R1_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R2_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R2_INV_1 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y22__R3_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B155));
  sky130_fd_sc_hd__clkbuf_4 T32Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2516));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R0_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2552));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R1_INV_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R2_INV_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R2_INV_1 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2588));
  sky130_fd_sc_hd__clkbuf_4 T32Y24__R0_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B164));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R0_INV_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2660));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R1_INV_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R2_INV_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R2_INV_1 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2696));
  sky130_fd_sc_hd__clkbuf_4 T32Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2732));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R0_INV_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y25__R1_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B173));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R1_INV_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R2_INV_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R2_INV_1 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2804));
  sky130_fd_sc_hd__clkbuf_4 T32Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2840));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R0_INV_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2876));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R1_INV_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R2_INV_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R2_INV_1 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y26__R3_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B182));
  sky130_fd_sc_hd__clkbuf_4 T32Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2948));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R0_INV_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2984));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R1_INV_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R2_INV_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R2_INV_1 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3020));
  sky130_fd_sc_hd__clkbuf_4 T32Y28__R0_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B191));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R0_INV_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3092));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R1_INV_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R2_INV_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R2_INV_1 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3128));
  sky130_fd_sc_hd__clkbuf_4 T32Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3164));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R0_INV_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y29__R1_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B200));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R1_INV_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R2_INV_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R2_INV_1 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3236));
  sky130_fd_sc_hd__clkbuf_4 T32Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B252));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R0_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y2__R1_BUF_0 (.A(clk_L1_B17), .X(clk_L0_B287));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R1_INV_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R2_INV_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R2_INV_1 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y2__R3_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B323));
  sky130_fd_sc_hd__clkbuf_4 T32Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3272));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R0_INV_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3308));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R1_INV_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R2_INV_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R2_INV_1 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y30__R3_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B209));
  sky130_fd_sc_hd__clkbuf_4 T32Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3380));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R0_INV_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3416));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R1_INV_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R2_INV_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R2_INV_1 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3452));
  sky130_fd_sc_hd__clkbuf_4 T32Y32__R0_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B218));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R0_INV_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3524));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R1_INV_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R2_INV_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R2_INV_1 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3560));
  sky130_fd_sc_hd__clkbuf_4 T32Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3596));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R0_INV_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y33__R1_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B227));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R1_INV_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R2_INV_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R2_INV_1 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3668));
  sky130_fd_sc_hd__clkbuf_4 T32Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3704));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R0_INV_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3740));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R1_INV_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R2_INV_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R2_INV_1 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y34__R3_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B236));
  sky130_fd_sc_hd__clkbuf_4 T32Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3812));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R0_INV_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3848));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R1_INV_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R2_INV_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R2_INV_1 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3884));
  sky130_fd_sc_hd__clkbuf_4 T32Y36__R0_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B245));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R0_INV_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3956));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R1_INV_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R2_INV_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R2_INV_1 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3992));
  sky130_fd_sc_hd__clkbuf_4 T32Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4028));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R0_INV_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y37__R1_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B254));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R1_INV_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R2_INV_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R2_INV_1 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4100));
  sky130_fd_sc_hd__clkbuf_4 T32Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4136));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R0_INV_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4172));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R1_INV_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R2_INV_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R2_INV_1 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y38__R3_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B263));
  sky130_fd_sc_hd__clkbuf_4 T32Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4244));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R0_INV_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4280));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R1_INV_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R2_INV_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R2_INV_1 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4316));
  sky130_fd_sc_hd__clkbuf_4 T32Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B358));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R0_INV_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B393));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R1_INV_0 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R2_INV_0 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R2_INV_1 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B429));
  sky130_fd_sc_hd__clkbuf_4 T32Y40__R0_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B17));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R0_INV_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4388));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R1_INV_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R2_INV_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R2_INV_1 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4424));
  sky130_fd_sc_hd__clkbuf_4 T32Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4460));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R0_INV_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y41__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B281));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R1_INV_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R2_INV_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R2_INV_1 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4532));
  sky130_fd_sc_hd__clkbuf_4 T32Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4568));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R0_INV_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4604));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R1_INV_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R2_INV_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R2_INV_1 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y42__R3_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B290));
  sky130_fd_sc_hd__clkbuf_4 T32Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4676));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R0_INV_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4712));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R1_INV_0 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R2_INV_0 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R2_INV_1 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4748));
  sky130_fd_sc_hd__clkbuf_4 T32Y44__R0_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B299));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R0_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4820));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R1_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R2_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R2_INV_1 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4856));
  sky130_fd_sc_hd__clkbuf_4 T32Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4892));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R0_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y45__R1_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B308));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R1_INV_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R2_INV_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R2_INV_1 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4964));
  sky130_fd_sc_hd__clkbuf_4 T32Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5000));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R0_INV_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5036));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R1_INV_0 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R2_INV_0 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R2_INV_1 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y46__R3_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B317));
  sky130_fd_sc_hd__clkbuf_4 T32Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5108));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R0_INV_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5144));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R1_INV_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R2_INV_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R2_INV_1 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5180));
  sky130_fd_sc_hd__clkbuf_4 T32Y48__R0_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B326));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R0_INV_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5252));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R1_INV_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R2_INV_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R2_INV_1 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5288));
  sky130_fd_sc_hd__clkbuf_4 T32Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5324));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R0_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y49__R1_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B335));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R1_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R2_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R2_INV_1 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5396));
  sky130_fd_sc_hd__clkbuf_4 T32Y4__R0_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B465));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R0_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B501));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R1_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R2_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R2_INV_1 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B537));
  sky130_fd_sc_hd__clkbuf_4 T32Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5432));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R0_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5468));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R1_INV_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R2_INV_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R2_INV_1 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y50__R3_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B344));
  sky130_fd_sc_hd__clkbuf_4 T32Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5540));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R0_INV_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5576));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R1_INV_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R2_INV_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R2_INV_1 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5612));
  sky130_fd_sc_hd__clkbuf_4 T32Y52__R0_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B353));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R0_INV_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5684));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R1_INV_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R2_INV_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R2_INV_1 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5720));
  sky130_fd_sc_hd__clkbuf_4 T32Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5756));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R0_INV_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y53__R1_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B362));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R1_INV_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R2_INV_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R2_INV_1 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5828));
  sky130_fd_sc_hd__clkbuf_4 T32Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5864));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R0_INV_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5900));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R1_INV_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R2_INV_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R2_INV_1 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y54__R3_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B371));
  sky130_fd_sc_hd__clkbuf_4 T32Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5972));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R0_INV_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6008));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R1_INV_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R2_INV_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R2_INV_1 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6044));
  sky130_fd_sc_hd__clkbuf_4 T32Y56__R0_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B380));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R0_INV_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6116));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R1_INV_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R2_INV_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R2_INV_1 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6152));
  sky130_fd_sc_hd__clkbuf_4 T32Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6188));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R0_INV_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y57__R1_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B389));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R1_INV_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R2_INV_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R2_INV_1 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6260));
  sky130_fd_sc_hd__clkbuf_4 T32Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6296));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R0_INV_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6332));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R1_INV_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R2_INV_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R2_INV_1 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y58__R3_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B398));
  sky130_fd_sc_hd__clkbuf_4 T32Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6404));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R0_INV_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6440));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R1_INV_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R2_INV_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R2_INV_1 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6476));
  sky130_fd_sc_hd__clkbuf_4 T32Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B573));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R0_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y5__R1_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B609));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R1_INV_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R2_INV_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R2_INV_1 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B645));
  sky130_fd_sc_hd__clkbuf_4 T32Y60__R0_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B407));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R0_INV_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6548));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R1_INV_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R2_INV_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R2_INV_1 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6584));
  sky130_fd_sc_hd__clkbuf_4 T32Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6620));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R0_INV_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y61__R1_BUF_0 (.A(clk_L4_B0), .X(clk_L3_B2));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R1_INV_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R2_INV_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R2_INV_1 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6692));
  sky130_fd_sc_hd__clkbuf_4 T32Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6728));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R0_INV_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6764));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R1_INV_0 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R2_INV_0 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R2_INV_1 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y62__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B425));
  sky130_fd_sc_hd__clkbuf_4 T32Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6836));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R0_INV_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6872));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R1_INV_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R2_INV_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R2_INV_1 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6908));
  sky130_fd_sc_hd__clkbuf_4 T32Y64__R0_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B434));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R0_INV_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6980));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R1_INV_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R2_INV_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R2_INV_1 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7016));
  sky130_fd_sc_hd__clkbuf_4 T32Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7052));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R0_INV_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y65__R1_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B443));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R1_INV_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R2_INV_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R2_INV_1 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7124));
  sky130_fd_sc_hd__clkbuf_4 T32Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7160));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R0_INV_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7196));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R1_INV_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R2_INV_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R2_INV_1 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y66__R3_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B452));
  sky130_fd_sc_hd__clkbuf_4 T32Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7268));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R0_INV_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7304));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R1_INV_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R2_INV_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R2_INV_1 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7340));
  sky130_fd_sc_hd__clkbuf_4 T32Y68__R0_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B461));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R0_INV_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7412));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R1_INV_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R2_INV_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R2_INV_1 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7448));
  sky130_fd_sc_hd__clkbuf_4 T32Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7484));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R0_INV_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y69__R1_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B470));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R1_INV_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R2_INV_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R2_INV_1 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7556));
  sky130_fd_sc_hd__clkbuf_4 T32Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B681));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R0_INV_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B717));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R1_INV_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R2_INV_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R2_INV_1 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y6__R3_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B753));
  sky130_fd_sc_hd__clkbuf_4 T32Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7592));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R0_INV_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7628));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R1_INV_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R2_INV_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R2_INV_1 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y70__R3_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B479));
  sky130_fd_sc_hd__clkbuf_4 T32Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7700));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R0_INV_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7736));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R1_INV_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R2_INV_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R2_INV_1 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7772));
  sky130_fd_sc_hd__clkbuf_4 T32Y72__R0_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B488));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R0_INV_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7844));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R1_INV_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R2_INV_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R2_INV_1 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7880));
  sky130_fd_sc_hd__clkbuf_4 T32Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7916));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R0_INV_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y73__R1_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B497));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R1_INV_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R2_INV_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R2_INV_1 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7988));
  sky130_fd_sc_hd__clkbuf_4 T32Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8024));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R0_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8060));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R1_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R2_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R2_INV_1 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y74__R3_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B506));
  sky130_fd_sc_hd__clkbuf_4 T32Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8132));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R0_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8168));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R1_INV_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R2_INV_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R2_INV_1 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8204));
  sky130_fd_sc_hd__clkbuf_4 T32Y76__R0_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B515));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R0_INV_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8276));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R1_INV_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R2_INV_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R2_INV_1 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8312));
  sky130_fd_sc_hd__clkbuf_4 T32Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8348));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R0_INV_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y77__R1_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B524));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R1_INV_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R2_INV_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R2_INV_1 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8420));
  sky130_fd_sc_hd__clkbuf_4 T32Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8456));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R0_INV_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8492));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R1_INV_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R2_INV_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R2_INV_1 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y78__R3_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B533));
  sky130_fd_sc_hd__clkbuf_4 T32Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8564));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R0_INV_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8600));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R1_INV_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R2_INV_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R2_INV_1 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8636));
  sky130_fd_sc_hd__clkbuf_4 T32Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B789));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R0_INV_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B825));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R1_INV_0 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R2_INV_0 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R2_INV_1 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B861));
  sky130_fd_sc_hd__clkbuf_4 T32Y80__R0_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B542));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R0_INV_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8708));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R1_INV_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R2_INV_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R2_INV_1 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8744));
  sky130_fd_sc_hd__clkbuf_4 T32Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8780));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R0_INV_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y81__R1_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B551));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R1_INV_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R2_INV_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R2_INV_1 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8852));
  sky130_fd_sc_hd__clkbuf_4 T32Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8888));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R0_INV_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8924));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R1_INV_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R2_INV_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R2_INV_1 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y82__R3_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B35));
  sky130_fd_sc_hd__clkbuf_4 T32Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8996));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R0_INV_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9032));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R1_INV_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R2_INV_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R2_INV_1 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9068));
  sky130_fd_sc_hd__clkbuf_4 T32Y84__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B569));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R0_INV_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9140));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R1_INV_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R2_INV_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R2_INV_1 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9176));
  sky130_fd_sc_hd__clkbuf_4 T32Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9212));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R0_INV_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y85__R1_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B578));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R1_INV_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R2_INV_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R2_INV_1 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9284));
  sky130_fd_sc_hd__clkbuf_4 T32Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9320));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R0_INV_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9356));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R1_INV_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R2_INV_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R2_INV_1 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y86__R3_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B587));
  sky130_fd_sc_hd__clkbuf_4 T32Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9428));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R0_INV_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9464));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R1_INV_0 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R2_INV_0 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R2_INV_1 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9500));
  sky130_fd_sc_hd__clkbuf_4 T32Y88__R0_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B596));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R0_INV_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9572));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R1_INV_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R2_INV_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R2_INV_1 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9608));
  sky130_fd_sc_hd__clkbuf_4 T32Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9644));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R0_INV_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y89__R1_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B605));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R1_INV_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R2_INV_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R2_INV_1 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9716));
  sky130_fd_sc_hd__clkbuf_4 T32Y8__R0_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B897));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R0_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B933));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R1_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R2_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R2_INV_1 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B969));
  sky130_fd_sc_hd__clkbuf_4 T32Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1005));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R0_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y9__R1_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1041));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R1_INV_0 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R2_INV_0 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R2_INV_1 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1077));
  sky130_fd_sc_hd__clkbuf_4 T33Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B43));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R0_INV_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B78));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R1_INV_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R2_INV_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R2_INV_1 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y0__R3_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B113));
  sky130_fd_sc_hd__clkbuf_4 T33Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1114));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R0_INV_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1150));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R1_INV_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R2_INV_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R2_INV_1 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y10__R3_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1186));
  sky130_fd_sc_hd__clkbuf_4 T33Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1222));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R0_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1258));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R1_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R2_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R2_INV_1 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1294));
  sky130_fd_sc_hd__clkbuf_4 T33Y12__R0_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1330));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R0_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1366));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R1_INV_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R2_INV_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R2_INV_1 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1402));
  sky130_fd_sc_hd__clkbuf_4 T33Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1438));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R0_INV_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y13__R1_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1474));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R1_INV_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R2_INV_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R2_INV_1 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1510));
  sky130_fd_sc_hd__clkbuf_4 T33Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1546));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R0_INV_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1581));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R1_INV_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R2_INV_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R2_INV_1 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y14__R3_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1617));
  sky130_fd_sc_hd__clkbuf_4 T33Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1653));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R0_INV_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1689));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R1_INV_0 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R2_INV_0 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R2_INV_1 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1725));
  sky130_fd_sc_hd__clkbuf_4 T33Y16__R0_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1761));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R0_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1797));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R1_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R2_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R2_INV_1 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1833));
  sky130_fd_sc_hd__clkbuf_4 T33Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1869));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R0_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y17__R1_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1905));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R1_INV_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R2_INV_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R2_INV_1 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1941));
  sky130_fd_sc_hd__clkbuf_4 T33Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1977));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R0_INV_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2013));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R1_INV_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R2_INV_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R2_INV_1 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y18__R3_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2049));
  sky130_fd_sc_hd__clkbuf_4 T33Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2085));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R0_INV_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2121));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R1_INV_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R2_INV_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R2_INV_1 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2157));
  sky130_fd_sc_hd__clkbuf_4 T33Y1__R0_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B148));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R0_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B183));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R1_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R2_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R2_INV_1 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B218));
  sky130_fd_sc_hd__clkbuf_4 T33Y20__R0_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2193));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R0_INV_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2229));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R1_INV_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R2_INV_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R2_INV_1 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2265));
  sky130_fd_sc_hd__clkbuf_4 T33Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2301));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R0_INV_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y21__R1_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2337));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R1_INV_0 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R2_INV_0 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R2_INV_1 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2373));
  sky130_fd_sc_hd__clkbuf_4 T33Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2409));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R0_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2445));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R1_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R2_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R2_INV_1 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y22__R3_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2481));
  sky130_fd_sc_hd__clkbuf_4 T33Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2517));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R0_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2553));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R1_INV_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R2_INV_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R2_INV_1 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2589));
  sky130_fd_sc_hd__clkbuf_4 T33Y24__R0_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2625));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R0_INV_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2661));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R1_INV_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R2_INV_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R2_INV_1 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2697));
  sky130_fd_sc_hd__clkbuf_4 T33Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2733));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R0_INV_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y25__R1_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2769));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R1_INV_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R2_INV_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R2_INV_1 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2805));
  sky130_fd_sc_hd__clkbuf_4 T33Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2841));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R0_INV_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2877));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R1_INV_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R2_INV_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R2_INV_1 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y26__R3_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2913));
  sky130_fd_sc_hd__clkbuf_4 T33Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2949));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R0_INV_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2985));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R1_INV_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R2_INV_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R2_INV_1 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3021));
  sky130_fd_sc_hd__clkbuf_4 T33Y28__R0_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3057));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R0_INV_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3093));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R1_INV_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R2_INV_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R2_INV_1 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3129));
  sky130_fd_sc_hd__clkbuf_4 T33Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3165));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R0_INV_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y29__R1_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3201));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R1_INV_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R2_INV_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R2_INV_1 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3237));
  sky130_fd_sc_hd__clkbuf_4 T33Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B253));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R0_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y2__R1_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B18));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R1_INV_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R2_INV_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R2_INV_1 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y2__R3_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B324));
  sky130_fd_sc_hd__clkbuf_4 T33Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3273));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R0_INV_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3309));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R1_INV_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R2_INV_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R2_INV_1 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y30__R3_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3345));
  sky130_fd_sc_hd__clkbuf_4 T33Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3381));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R0_INV_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3417));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R1_INV_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R2_INV_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R2_INV_1 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3453));
  sky130_fd_sc_hd__clkbuf_4 T33Y32__R0_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3489));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R0_INV_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3525));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R1_INV_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R2_INV_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R2_INV_1 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3561));
  sky130_fd_sc_hd__clkbuf_4 T33Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3597));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R0_INV_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y33__R1_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3633));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R1_INV_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R2_INV_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R2_INV_1 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3669));
  sky130_fd_sc_hd__clkbuf_4 T33Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3705));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R0_INV_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3741));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R1_INV_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R2_INV_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R2_INV_1 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y34__R3_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3777));
  sky130_fd_sc_hd__clkbuf_4 T33Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3813));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R0_INV_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3849));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R1_INV_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R2_INV_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R2_INV_1 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3885));
  sky130_fd_sc_hd__clkbuf_4 T33Y36__R0_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3921));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R0_INV_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3957));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R1_INV_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R2_INV_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R2_INV_1 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3993));
  sky130_fd_sc_hd__clkbuf_4 T33Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4029));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R0_INV_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y37__R1_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4065));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R1_INV_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R2_INV_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R2_INV_1 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4101));
  sky130_fd_sc_hd__clkbuf_4 T33Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4137));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R0_INV_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4173));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R1_INV_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R2_INV_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R2_INV_1 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y38__R3_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4209));
  sky130_fd_sc_hd__clkbuf_4 T33Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4245));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R0_INV_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4281));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R1_INV_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R2_INV_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R2_INV_1 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4317));
  sky130_fd_sc_hd__clkbuf_4 T33Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B359));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R0_INV_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B394));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R1_INV_0 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R2_INV_0 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R2_INV_1 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B430));
  sky130_fd_sc_hd__clkbuf_4 T33Y40__R0_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4353));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R0_INV_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4389));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R1_INV_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R2_INV_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R2_INV_1 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4425));
  sky130_fd_sc_hd__clkbuf_4 T33Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4461));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R0_INV_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y41__R1_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4497));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R1_INV_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R2_INV_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R2_INV_1 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4533));
  sky130_fd_sc_hd__clkbuf_4 T33Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4569));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R0_INV_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4605));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R1_INV_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R2_INV_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R2_INV_1 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y42__R3_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4641));
  sky130_fd_sc_hd__clkbuf_4 T33Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4677));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R0_INV_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4713));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R1_INV_0 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R2_INV_0 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R2_INV_1 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4749));
  sky130_fd_sc_hd__clkbuf_4 T33Y44__R0_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4785));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R0_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4821));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R1_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R2_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R2_INV_1 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4857));
  sky130_fd_sc_hd__clkbuf_4 T33Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4893));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R0_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y45__R1_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4929));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R1_INV_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R2_INV_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R2_INV_1 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4965));
  sky130_fd_sc_hd__clkbuf_4 T33Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5001));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R0_INV_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5037));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R1_INV_0 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R2_INV_0 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R2_INV_1 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y46__R3_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5073));
  sky130_fd_sc_hd__clkbuf_4 T33Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5109));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R0_INV_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5145));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R1_INV_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R2_INV_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R2_INV_1 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5181));
  sky130_fd_sc_hd__clkbuf_4 T33Y48__R0_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5217));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R0_INV_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5253));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R1_INV_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R2_INV_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R2_INV_1 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5289));
  sky130_fd_sc_hd__clkbuf_4 T33Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5325));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R0_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y49__R1_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5361));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R1_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R2_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R2_INV_1 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5397));
  sky130_fd_sc_hd__clkbuf_4 T33Y4__R0_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B466));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R0_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B502));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R1_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R2_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R2_INV_1 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B538));
  sky130_fd_sc_hd__clkbuf_4 T33Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5433));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R0_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5469));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R1_INV_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R2_INV_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R2_INV_1 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y50__R3_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5505));
  sky130_fd_sc_hd__clkbuf_4 T33Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5541));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R0_INV_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5577));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R1_INV_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R2_INV_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R2_INV_1 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5613));
  sky130_fd_sc_hd__clkbuf_4 T33Y52__R0_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5649));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R0_INV_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5685));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R1_INV_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R2_INV_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R2_INV_1 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5721));
  sky130_fd_sc_hd__clkbuf_4 T33Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5757));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R0_INV_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y53__R1_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5793));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R1_INV_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R2_INV_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R2_INV_1 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5829));
  sky130_fd_sc_hd__clkbuf_4 T33Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5865));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R0_INV_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5901));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R1_INV_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R2_INV_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R2_INV_1 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y54__R3_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5937));
  sky130_fd_sc_hd__clkbuf_4 T33Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5973));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R0_INV_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6009));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R1_INV_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R2_INV_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R2_INV_1 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6045));
  sky130_fd_sc_hd__clkbuf_4 T33Y56__R0_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6081));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R0_INV_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6117));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R1_INV_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R2_INV_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R2_INV_1 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6153));
  sky130_fd_sc_hd__clkbuf_4 T33Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6189));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R0_INV_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y57__R1_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6225));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R1_INV_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R2_INV_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R2_INV_1 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6261));
  sky130_fd_sc_hd__clkbuf_4 T33Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6297));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R0_INV_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6333));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R1_INV_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R2_INV_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R2_INV_1 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y58__R3_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6369));
  sky130_fd_sc_hd__clkbuf_4 T33Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6405));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R0_INV_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6441));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R1_INV_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R2_INV_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R2_INV_1 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6477));
  sky130_fd_sc_hd__clkbuf_4 T33Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B574));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R0_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y5__R1_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B610));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R1_INV_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R2_INV_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R2_INV_1 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B646));
  sky130_fd_sc_hd__clkbuf_4 T33Y60__R0_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6513));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R0_INV_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6549));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R1_INV_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R2_INV_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R2_INV_1 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6585));
  sky130_fd_sc_hd__clkbuf_4 T33Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6621));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R0_INV_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y61__R1_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6657));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R1_INV_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R2_INV_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R2_INV_1 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6693));
  sky130_fd_sc_hd__clkbuf_4 T33Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6729));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R0_INV_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6765));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R1_INV_0 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R2_INV_0 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R2_INV_1 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y62__R3_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6801));
  sky130_fd_sc_hd__clkbuf_4 T33Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6837));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R0_INV_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6873));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R1_INV_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R2_INV_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R2_INV_1 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6909));
  sky130_fd_sc_hd__clkbuf_4 T33Y64__R0_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6945));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R0_INV_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6981));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R1_INV_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R2_INV_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R2_INV_1 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7017));
  sky130_fd_sc_hd__clkbuf_4 T33Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7053));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R0_INV_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y65__R1_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7089));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R1_INV_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R2_INV_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R2_INV_1 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7125));
  sky130_fd_sc_hd__clkbuf_4 T33Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7161));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R0_INV_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7197));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R1_INV_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R2_INV_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R2_INV_1 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y66__R3_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7233));
  sky130_fd_sc_hd__clkbuf_4 T33Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7269));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R0_INV_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7305));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R1_INV_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R2_INV_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R2_INV_1 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7341));
  sky130_fd_sc_hd__clkbuf_4 T33Y68__R0_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7377));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R0_INV_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7413));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R1_INV_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R2_INV_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R2_INV_1 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7449));
  sky130_fd_sc_hd__clkbuf_4 T33Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7485));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R0_INV_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y69__R1_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7521));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R1_INV_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R2_INV_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R2_INV_1 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7557));
  sky130_fd_sc_hd__clkbuf_4 T33Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B682));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R0_INV_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B718));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R1_INV_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R2_INV_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R2_INV_1 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y6__R3_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B754));
  sky130_fd_sc_hd__clkbuf_4 T33Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7593));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R0_INV_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7629));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R1_INV_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R2_INV_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R2_INV_1 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y70__R3_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7665));
  sky130_fd_sc_hd__clkbuf_4 T33Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7701));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R0_INV_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7737));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R1_INV_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R2_INV_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R2_INV_1 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7773));
  sky130_fd_sc_hd__clkbuf_4 T33Y72__R0_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7809));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R0_INV_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7845));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R1_INV_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R2_INV_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R2_INV_1 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7881));
  sky130_fd_sc_hd__clkbuf_4 T33Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7917));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R0_INV_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y73__R1_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7953));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R1_INV_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R2_INV_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R2_INV_1 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7989));
  sky130_fd_sc_hd__clkbuf_4 T33Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8025));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R0_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8061));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R1_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R2_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R2_INV_1 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y74__R3_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8097));
  sky130_fd_sc_hd__clkbuf_4 T33Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8133));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R0_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8169));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R1_INV_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R2_INV_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R2_INV_1 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8205));
  sky130_fd_sc_hd__clkbuf_4 T33Y76__R0_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8241));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R0_INV_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8277));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R1_INV_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R2_INV_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R2_INV_1 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8313));
  sky130_fd_sc_hd__clkbuf_4 T33Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8349));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R0_INV_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y77__R1_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8385));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R1_INV_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R2_INV_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R2_INV_1 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8421));
  sky130_fd_sc_hd__clkbuf_4 T33Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8457));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R0_INV_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8493));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R1_INV_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R2_INV_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R2_INV_1 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y78__R3_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8529));
  sky130_fd_sc_hd__clkbuf_4 T33Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8565));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R0_INV_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8601));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R1_INV_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R2_INV_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R2_INV_1 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8637));
  sky130_fd_sc_hd__clkbuf_4 T33Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B790));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R0_INV_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B826));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R1_INV_0 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R2_INV_0 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R2_INV_1 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B862));
  sky130_fd_sc_hd__clkbuf_4 T33Y80__R0_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8673));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R0_INV_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8709));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R1_INV_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R2_INV_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R2_INV_1 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8745));
  sky130_fd_sc_hd__clkbuf_4 T33Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8781));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R0_INV_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y81__R1_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8817));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R1_INV_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R2_INV_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R2_INV_1 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8853));
  sky130_fd_sc_hd__clkbuf_4 T33Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8889));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R0_INV_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8925));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R1_INV_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R2_INV_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R2_INV_1 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y82__R3_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8961));
  sky130_fd_sc_hd__clkbuf_4 T33Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8997));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R0_INV_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9033));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R1_INV_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R2_INV_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R2_INV_1 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9069));
  sky130_fd_sc_hd__clkbuf_4 T33Y84__R0_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9105));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R0_INV_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9141));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R1_INV_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R2_INV_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R2_INV_1 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9177));
  sky130_fd_sc_hd__clkbuf_4 T33Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9213));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R0_INV_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y85__R1_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9249));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R1_INV_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R2_INV_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R2_INV_1 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9285));
  sky130_fd_sc_hd__clkbuf_4 T33Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9321));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R0_INV_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9357));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R1_INV_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R2_INV_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R2_INV_1 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y86__R3_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9393));
  sky130_fd_sc_hd__clkbuf_4 T33Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9429));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R0_INV_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9465));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R1_INV_0 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R2_INV_0 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R2_INV_1 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9501));
  sky130_fd_sc_hd__clkbuf_4 T33Y88__R0_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9537));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R0_INV_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9573));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R1_INV_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R2_INV_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R2_INV_1 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9609));
  sky130_fd_sc_hd__clkbuf_4 T33Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9645));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R0_INV_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y89__R1_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9681));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R1_INV_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R2_INV_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R2_INV_1 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9717));
  sky130_fd_sc_hd__clkbuf_4 T33Y8__R0_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B898));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R0_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B934));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R1_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R2_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R2_INV_1 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B970));
  sky130_fd_sc_hd__clkbuf_4 T33Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1006));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R0_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y9__R1_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1042));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R1_INV_0 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R2_INV_0 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R2_INV_1 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1078));
  sky130_fd_sc_hd__clkbuf_4 T34Y0__R0_BUF_0 (.A(clk_L1_B2), .X(clk_L0_B44));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R0_INV_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y0__R1_BUF_0 (.A(clk_L1_B4), .X(clk_L0_B79));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R1_INV_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R2_INV_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R2_INV_1 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y0__R3_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B114));
  sky130_fd_sc_hd__clkbuf_4 T34Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1115));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R0_INV_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y10__R1_BUF_0 (.A(clk_L1_B71), .X(clk_L0_B1151));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R1_INV_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R2_INV_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R2_INV_1 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y10__R3_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1187));
  sky130_fd_sc_hd__clkbuf_4 T34Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1223));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R0_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1259));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R1_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R2_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R2_INV_1 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y11__R3_BUF_0 (.A(clk_L1_B80), .X(clk_L0_B1295));
  sky130_fd_sc_hd__clkbuf_4 T34Y12__R0_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1331));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R0_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1367));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R1_INV_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R2_INV_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R2_INV_1 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1403));
  sky130_fd_sc_hd__clkbuf_4 T34Y13__R0_BUF_0 (.A(clk_L1_B89), .X(clk_L0_B1439));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R0_INV_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y13__R1_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1475));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R1_INV_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R2_INV_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R2_INV_1 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1511));
  sky130_fd_sc_hd__clkbuf_4 T34Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1547));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R0_INV_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1582));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R1_INV_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R2_INV_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R2_INV_1 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y14__R3_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1618));
  sky130_fd_sc_hd__clkbuf_4 T34Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1654));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R0_INV_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1690));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R1_INV_0 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R2_INV_0 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R2_INV_1 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1726));
  sky130_fd_sc_hd__clkbuf_4 T34Y16__R0_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1762));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R0_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1798));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R1_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R2_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R2_INV_1 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1834));
  sky130_fd_sc_hd__clkbuf_4 T34Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1870));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R0_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y17__R1_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1906));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R1_INV_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R2_INV_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R2_INV_1 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1942));
  sky130_fd_sc_hd__clkbuf_4 T34Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1978));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R0_INV_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2014));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R1_INV_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R2_INV_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R2_INV_1 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y18__R3_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2050));
  sky130_fd_sc_hd__clkbuf_4 T34Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2086));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R0_INV_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2122));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R1_INV_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R2_INV_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R2_INV_1 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2158));
  sky130_fd_sc_hd__clkbuf_4 T34Y1__R0_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B149));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R0_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y1__R1_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B184));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R1_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R2_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R2_INV_1 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y1__R3_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B219));
  sky130_fd_sc_hd__clkbuf_4 T34Y20__R0_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2194));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R0_INV_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2230));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R1_INV_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R2_INV_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R2_INV_1 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2266));
  sky130_fd_sc_hd__clkbuf_4 T34Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2302));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R0_INV_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y21__R1_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2338));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R1_INV_0 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R2_INV_0 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R2_INV_1 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2374));
  sky130_fd_sc_hd__clkbuf_4 T34Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2410));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R0_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2446));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R1_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R2_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R2_INV_1 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y22__R3_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2482));
  sky130_fd_sc_hd__clkbuf_4 T34Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2518));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R0_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2554));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R1_INV_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R2_INV_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R2_INV_1 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2590));
  sky130_fd_sc_hd__clkbuf_4 T34Y24__R0_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2626));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R0_INV_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2662));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R1_INV_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R2_INV_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R2_INV_1 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2698));
  sky130_fd_sc_hd__clkbuf_4 T34Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2734));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R0_INV_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y25__R1_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2770));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R1_INV_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R2_INV_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R2_INV_1 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2806));
  sky130_fd_sc_hd__clkbuf_4 T34Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2842));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R0_INV_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2878));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R1_INV_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R2_INV_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R2_INV_1 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y26__R3_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2914));
  sky130_fd_sc_hd__clkbuf_4 T34Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2950));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R0_INV_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2986));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R1_INV_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R2_INV_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R2_INV_1 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3022));
  sky130_fd_sc_hd__clkbuf_4 T34Y28__R0_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3058));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R0_INV_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3094));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R1_INV_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R2_INV_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R2_INV_1 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3130));
  sky130_fd_sc_hd__clkbuf_4 T34Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3166));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R0_INV_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y29__R1_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3202));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R1_INV_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R2_INV_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R2_INV_1 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3238));
  sky130_fd_sc_hd__clkbuf_4 T34Y2__R0_BUF_0 (.A(clk_L1_B15), .X(clk_L0_B254));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R0_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y2__R1_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B289));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R1_INV_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R2_INV_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R2_INV_1 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y2__R3_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B325));
  sky130_fd_sc_hd__clkbuf_4 T34Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3274));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R0_INV_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3310));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R1_INV_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R2_INV_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R2_INV_1 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y30__R3_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3346));
  sky130_fd_sc_hd__clkbuf_4 T34Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3382));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R0_INV_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3418));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R1_INV_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R2_INV_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R2_INV_1 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3454));
  sky130_fd_sc_hd__clkbuf_4 T34Y32__R0_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3490));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R0_INV_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3526));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R1_INV_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R2_INV_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R2_INV_1 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3562));
  sky130_fd_sc_hd__clkbuf_4 T34Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3598));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R0_INV_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y33__R1_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3634));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R1_INV_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R2_INV_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R2_INV_1 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3670));
  sky130_fd_sc_hd__clkbuf_4 T34Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3706));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R0_INV_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3742));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R1_INV_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R2_INV_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R2_INV_1 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y34__R3_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3778));
  sky130_fd_sc_hd__clkbuf_4 T34Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3814));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R0_INV_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3850));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R1_INV_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R2_INV_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R2_INV_1 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3886));
  sky130_fd_sc_hd__clkbuf_4 T34Y36__R0_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3922));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R0_INV_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3958));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R1_INV_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R2_INV_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R2_INV_1 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3994));
  sky130_fd_sc_hd__clkbuf_4 T34Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4030));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R0_INV_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y37__R1_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4066));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R1_INV_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R2_INV_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R2_INV_1 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4102));
  sky130_fd_sc_hd__clkbuf_4 T34Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4138));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R0_INV_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4174));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R1_INV_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R2_INV_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R2_INV_1 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y38__R3_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4210));
  sky130_fd_sc_hd__clkbuf_4 T34Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4246));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R0_INV_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4282));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R1_INV_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R2_INV_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R2_INV_1 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4318));
  sky130_fd_sc_hd__clkbuf_4 T34Y3__R0_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B360));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R0_INV_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B395));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R1_INV_0 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R2_INV_0 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R2_INV_1 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y3__R3_BUF_0 (.A(clk_L1_B26), .X(clk_L0_B431));
  sky130_fd_sc_hd__clkbuf_4 T34Y40__R0_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4354));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R0_INV_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4390));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R1_INV_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R2_INV_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R2_INV_1 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4426));
  sky130_fd_sc_hd__clkbuf_4 T34Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4462));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R0_INV_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y41__R1_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4498));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R1_INV_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R2_INV_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R2_INV_1 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4534));
  sky130_fd_sc_hd__clkbuf_4 T34Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4570));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R0_INV_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4606));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R1_INV_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R2_INV_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R2_INV_1 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y42__R3_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4642));
  sky130_fd_sc_hd__clkbuf_4 T34Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4678));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R0_INV_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4714));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R1_INV_0 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R2_INV_0 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R2_INV_1 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4750));
  sky130_fd_sc_hd__clkbuf_4 T34Y44__R0_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4786));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R0_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4822));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R1_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R2_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R2_INV_1 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4858));
  sky130_fd_sc_hd__clkbuf_4 T34Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4894));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R0_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y45__R1_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4930));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R1_INV_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R2_INV_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R2_INV_1 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4966));
  sky130_fd_sc_hd__clkbuf_4 T34Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5002));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R0_INV_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5038));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R1_INV_0 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R2_INV_0 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R2_INV_1 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y46__R3_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5074));
  sky130_fd_sc_hd__clkbuf_4 T34Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5110));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R0_INV_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5146));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R1_INV_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R2_INV_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R2_INV_1 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5182));
  sky130_fd_sc_hd__clkbuf_4 T34Y48__R0_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5218));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R0_INV_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5254));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R1_INV_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R2_INV_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R2_INV_1 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5290));
  sky130_fd_sc_hd__clkbuf_4 T34Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5326));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R0_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y49__R1_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5362));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R1_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R2_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R2_INV_1 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5398));
  sky130_fd_sc_hd__clkbuf_4 T34Y4__R0_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B467));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R0_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B503));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R1_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R2_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R2_INV_1 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B539));
  sky130_fd_sc_hd__clkbuf_4 T34Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5434));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R0_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5470));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R1_INV_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R2_INV_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R2_INV_1 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y50__R3_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5506));
  sky130_fd_sc_hd__clkbuf_4 T34Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5542));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R0_INV_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5578));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R1_INV_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R2_INV_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R2_INV_1 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5614));
  sky130_fd_sc_hd__clkbuf_4 T34Y52__R0_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5650));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R0_INV_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5686));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R1_INV_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R2_INV_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R2_INV_1 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5722));
  sky130_fd_sc_hd__clkbuf_4 T34Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5758));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R0_INV_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y53__R1_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5794));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R1_INV_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R2_INV_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R2_INV_1 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5830));
  sky130_fd_sc_hd__clkbuf_4 T34Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5866));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R0_INV_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5902));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R1_INV_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R2_INV_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R2_INV_1 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y54__R3_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5938));
  sky130_fd_sc_hd__clkbuf_4 T34Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5974));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R0_INV_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6010));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R1_INV_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R2_INV_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R2_INV_1 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6046));
  sky130_fd_sc_hd__clkbuf_4 T34Y56__R0_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6082));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R0_INV_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6118));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R1_INV_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R2_INV_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R2_INV_1 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6154));
  sky130_fd_sc_hd__clkbuf_4 T34Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6190));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R0_INV_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y57__R1_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6226));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R1_INV_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R2_INV_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R2_INV_1 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6262));
  sky130_fd_sc_hd__clkbuf_4 T34Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6298));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R0_INV_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6334));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R1_INV_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R2_INV_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R2_INV_1 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y58__R3_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6370));
  sky130_fd_sc_hd__clkbuf_4 T34Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6406));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R0_INV_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6442));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R1_INV_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R2_INV_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R2_INV_1 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6478));
  sky130_fd_sc_hd__clkbuf_4 T34Y5__R0_BUF_0 (.A(clk_L1_B35), .X(clk_L0_B575));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R0_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y5__R1_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B611));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R1_INV_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R2_INV_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R2_INV_1 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B647));
  sky130_fd_sc_hd__clkbuf_4 T34Y60__R0_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6514));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R0_INV_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6550));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R1_INV_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R2_INV_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R2_INV_1 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6586));
  sky130_fd_sc_hd__clkbuf_4 T34Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6622));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R0_INV_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y61__R1_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6658));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R1_INV_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R2_INV_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R2_INV_1 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6694));
  sky130_fd_sc_hd__clkbuf_4 T34Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6730));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R0_INV_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6766));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R1_INV_0 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R2_INV_0 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R2_INV_1 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y62__R3_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6802));
  sky130_fd_sc_hd__clkbuf_4 T34Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6838));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R0_INV_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6874));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R1_INV_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R2_INV_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R2_INV_1 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6910));
  sky130_fd_sc_hd__clkbuf_4 T34Y64__R0_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6946));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R0_INV_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6982));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R1_INV_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R2_INV_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R2_INV_1 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7018));
  sky130_fd_sc_hd__clkbuf_4 T34Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7054));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R0_INV_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y65__R1_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7090));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R1_INV_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R2_INV_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R2_INV_1 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7126));
  sky130_fd_sc_hd__clkbuf_4 T34Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7162));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R0_INV_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7198));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R1_INV_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R2_INV_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R2_INV_1 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y66__R3_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7234));
  sky130_fd_sc_hd__clkbuf_4 T34Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7270));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R0_INV_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7306));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R1_INV_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R2_INV_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R2_INV_1 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7342));
  sky130_fd_sc_hd__clkbuf_4 T34Y68__R0_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7378));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R0_INV_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7414));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R1_INV_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R2_INV_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R2_INV_1 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7450));
  sky130_fd_sc_hd__clkbuf_4 T34Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7486));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R0_INV_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y69__R1_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7522));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R1_INV_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R2_INV_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R2_INV_1 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7558));
  sky130_fd_sc_hd__clkbuf_4 T34Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B683));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R0_INV_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y6__R1_BUF_0 (.A(clk_L1_B44), .X(clk_L0_B719));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R1_INV_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R2_INV_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R2_INV_1 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y6__R3_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B755));
  sky130_fd_sc_hd__clkbuf_4 T34Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7594));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R0_INV_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7630));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R1_INV_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R2_INV_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R2_INV_1 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y70__R3_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7666));
  sky130_fd_sc_hd__clkbuf_4 T34Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7702));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R0_INV_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7738));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R1_INV_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R2_INV_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R2_INV_1 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7774));
  sky130_fd_sc_hd__clkbuf_4 T34Y72__R0_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7810));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R0_INV_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7846));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R1_INV_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R2_INV_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R2_INV_1 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7882));
  sky130_fd_sc_hd__clkbuf_4 T34Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7918));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R0_INV_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y73__R1_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7954));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R1_INV_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R2_INV_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R2_INV_1 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7990));
  sky130_fd_sc_hd__clkbuf_4 T34Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8026));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R0_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8062));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R1_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R2_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R2_INV_1 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y74__R3_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8098));
  sky130_fd_sc_hd__clkbuf_4 T34Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8134));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R0_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8170));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R1_INV_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R2_INV_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R2_INV_1 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8206));
  sky130_fd_sc_hd__clkbuf_4 T34Y76__R0_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8242));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R0_INV_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8278));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R1_INV_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R2_INV_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R2_INV_1 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8314));
  sky130_fd_sc_hd__clkbuf_4 T34Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8350));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R0_INV_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y77__R1_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8386));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R1_INV_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R2_INV_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R2_INV_1 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8422));
  sky130_fd_sc_hd__clkbuf_4 T34Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8458));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R0_INV_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8494));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R1_INV_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R2_INV_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R2_INV_1 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y78__R3_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8530));
  sky130_fd_sc_hd__clkbuf_4 T34Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8566));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R0_INV_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8602));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R1_INV_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R2_INV_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R2_INV_1 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8638));
  sky130_fd_sc_hd__clkbuf_4 T34Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B791));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R0_INV_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B827));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R1_INV_0 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R2_INV_0 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R2_INV_1 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y7__R3_BUF_0 (.A(clk_L1_B53), .X(clk_L0_B863));
  sky130_fd_sc_hd__clkbuf_4 T34Y80__R0_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8674));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R0_INV_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8710));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R1_INV_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R2_INV_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R2_INV_1 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8746));
  sky130_fd_sc_hd__clkbuf_4 T34Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8782));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R0_INV_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y81__R1_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8818));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R1_INV_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R2_INV_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R2_INV_1 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8854));
  sky130_fd_sc_hd__clkbuf_4 T34Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8890));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R0_INV_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8926));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R1_INV_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R2_INV_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R2_INV_1 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y82__R3_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8962));
  sky130_fd_sc_hd__clkbuf_4 T34Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8998));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R0_INV_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9034));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R1_INV_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R2_INV_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R2_INV_1 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9070));
  sky130_fd_sc_hd__clkbuf_4 T34Y84__R0_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9106));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R0_INV_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9142));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R1_INV_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R2_INV_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R2_INV_1 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9178));
  sky130_fd_sc_hd__clkbuf_4 T34Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9214));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R0_INV_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y85__R1_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9250));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R1_INV_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R2_INV_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R2_INV_1 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9286));
  sky130_fd_sc_hd__clkbuf_4 T34Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9322));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R0_INV_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9358));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R1_INV_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R2_INV_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R2_INV_1 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y86__R3_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9394));
  sky130_fd_sc_hd__clkbuf_4 T34Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9430));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R0_INV_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9466));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R1_INV_0 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R2_INV_0 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R2_INV_1 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9502));
  sky130_fd_sc_hd__clkbuf_4 T34Y88__R0_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9538));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R0_INV_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9574));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R1_INV_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R2_INV_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R2_INV_1 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9610));
  sky130_fd_sc_hd__clkbuf_4 T34Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9646));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R0_INV_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y89__R1_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9682));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R1_INV_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R2_INV_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R2_INV_1 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9718));
  sky130_fd_sc_hd__clkbuf_4 T34Y8__R0_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B899));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R0_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B935));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R1_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R2_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R2_INV_1 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B971));
  sky130_fd_sc_hd__clkbuf_4 T34Y9__R0_BUF_0 (.A(clk_L1_B62), .X(clk_L0_B1007));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R0_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y9__R1_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1043));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R1_INV_0 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R2_INV_0 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R2_INV_1 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1079));
  sky130_fd_sc_hd__clkbuf_4 T35Y0__R0_BUF_0 (.A(clk), .X(clk_L4_B0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R0_INV_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y0__R1_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B6));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R1_INV_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R2_INV_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R2_INV_1 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y0__R3_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B1));
  sky130_fd_sc_hd__clkbuf_4 T35Y10__R0_BUF_0 (.A(clk_L1_B69), .X(clk_L0_B1116));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R0_INV_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y10__R1_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B72));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R1_INV_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R2_INV_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R2_INV_1 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y10__R3_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1188));
  sky130_fd_sc_hd__clkbuf_4 T35Y11__R0_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1224));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R0_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y11__R1_BUF_0 (.A(clk_L1_B78), .X(clk_L0_B1260));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R1_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R2_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R2_INV_1 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y11__R3_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B81));
  sky130_fd_sc_hd__clkbuf_4 T35Y12__R0_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1332));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R0_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y12__R1_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1368));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R1_INV_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R2_INV_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R2_INV_1 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y12__R3_BUF_0 (.A(clk_L1_B87), .X(clk_L0_B1404));
  sky130_fd_sc_hd__clkbuf_4 T35Y13__R0_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B90));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R0_INV_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y13__R1_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1476));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R1_INV_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R2_INV_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R2_INV_1 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y13__R3_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1512));
  sky130_fd_sc_hd__clkbuf_4 T35Y14__R0_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1548));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R0_INV_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y14__R1_BUF_0 (.A(clk_L1_B98), .X(clk_L0_B1583));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R1_INV_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R2_INV_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R2_INV_1 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y14__R3_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1619));
  sky130_fd_sc_hd__clkbuf_4 T35Y15__R0_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1655));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R0_INV_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y15__R1_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1691));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R1_INV_0 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R2_INV_0 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R2_INV_1 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y15__R3_BUF_0 (.A(clk_L1_B107), .X(clk_L0_B1727));
  sky130_fd_sc_hd__clkbuf_4 T35Y16__R0_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1763));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R0_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y16__R1_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1799));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R1_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R2_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R2_INV_1 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y16__R3_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1835));
  sky130_fd_sc_hd__clkbuf_4 T35Y17__R0_BUF_0 (.A(clk_L1_B116), .X(clk_L0_B1871));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R0_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y17__R1_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1907));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R1_INV_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R2_INV_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R2_INV_1 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y17__R3_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1943));
  sky130_fd_sc_hd__clkbuf_4 T35Y18__R0_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1979));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R0_INV_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y18__R1_BUF_0 (.A(clk_L1_B125), .X(clk_L0_B2015));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R1_INV_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R2_INV_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R2_INV_1 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y18__R3_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2051));
  sky130_fd_sc_hd__clkbuf_4 T35Y19__R0_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2087));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R0_INV_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y19__R1_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2123));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R1_INV_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R2_INV_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R2_INV_1 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y19__R3_BUF_0 (.A(clk_L1_B134), .X(clk_L0_B2159));
  sky130_fd_sc_hd__clkbuf_4 T35Y1__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B2));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R0_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y1__R1_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B7));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R1_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R2_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R2_INV_1 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y1__R3_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B4));
  sky130_fd_sc_hd__clkbuf_4 T35Y20__R0_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2195));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R0_INV_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y20__R1_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2231));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R1_INV_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R2_INV_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R2_INV_1 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y20__R3_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2267));
  sky130_fd_sc_hd__clkbuf_4 T35Y21__R0_BUF_0 (.A(clk_L1_B143), .X(clk_L0_B2303));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R0_INV_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y21__R1_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2339));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R1_INV_0 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R2_INV_0 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R2_INV_1 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y21__R3_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2375));
  sky130_fd_sc_hd__clkbuf_4 T35Y22__R0_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2411));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R0_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y22__R1_BUF_0 (.A(clk_L1_B152), .X(clk_L0_B2447));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R1_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R2_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R2_INV_1 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y22__R3_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2483));
  sky130_fd_sc_hd__clkbuf_4 T35Y23__R0_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2519));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R0_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y23__R1_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2555));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R1_INV_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R2_INV_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R2_INV_1 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y23__R3_BUF_0 (.A(clk_L1_B161), .X(clk_L0_B2591));
  sky130_fd_sc_hd__clkbuf_4 T35Y24__R0_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2627));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R0_INV_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y24__R1_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2663));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R1_INV_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R2_INV_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R2_INV_1 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y24__R3_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2699));
  sky130_fd_sc_hd__clkbuf_4 T35Y25__R0_BUF_0 (.A(clk_L1_B170), .X(clk_L0_B2735));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R0_INV_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y25__R1_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2771));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R1_INV_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R2_INV_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R2_INV_1 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y25__R3_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2807));
  sky130_fd_sc_hd__clkbuf_4 T35Y26__R0_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2843));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R0_INV_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y26__R1_BUF_0 (.A(clk_L1_B179), .X(clk_L0_B2879));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R1_INV_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R2_INV_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R2_INV_1 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y26__R3_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2915));
  sky130_fd_sc_hd__clkbuf_4 T35Y27__R0_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2951));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R0_INV_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y27__R1_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2987));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R1_INV_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R2_INV_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R2_INV_1 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y27__R3_BUF_0 (.A(clk_L1_B188), .X(clk_L0_B3023));
  sky130_fd_sc_hd__clkbuf_4 T35Y28__R0_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3059));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R0_INV_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y28__R1_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3095));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R1_INV_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R2_INV_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R2_INV_1 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y28__R3_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3131));
  sky130_fd_sc_hd__clkbuf_4 T35Y29__R0_BUF_0 (.A(clk_L1_B197), .X(clk_L0_B3167));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R0_INV_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y29__R1_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3203));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R1_INV_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R2_INV_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R2_INV_1 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y29__R3_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3239));
  sky130_fd_sc_hd__clkbuf_4 T35Y2__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B5));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R0_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y2__R1_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B290));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R1_INV_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R2_INV_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R2_INV_1 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y2__R3_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B8));
  sky130_fd_sc_hd__clkbuf_4 T35Y30__R0_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3275));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R0_INV_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y30__R1_BUF_0 (.A(clk_L1_B206), .X(clk_L0_B3311));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R1_INV_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R2_INV_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R2_INV_1 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y30__R3_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3347));
  sky130_fd_sc_hd__clkbuf_4 T35Y31__R0_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3383));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R0_INV_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y31__R1_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3419));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R1_INV_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R2_INV_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R2_INV_1 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y31__R3_BUF_0 (.A(clk_L1_B215), .X(clk_L0_B3455));
  sky130_fd_sc_hd__clkbuf_4 T35Y32__R0_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3491));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R0_INV_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y32__R1_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3527));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R1_INV_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R2_INV_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R2_INV_1 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y32__R3_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3563));
  sky130_fd_sc_hd__clkbuf_4 T35Y33__R0_BUF_0 (.A(clk_L1_B224), .X(clk_L0_B3599));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R0_INV_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y33__R1_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3635));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R1_INV_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R2_INV_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R2_INV_1 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y33__R3_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3671));
  sky130_fd_sc_hd__clkbuf_4 T35Y34__R0_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3707));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R0_INV_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y34__R1_BUF_0 (.A(clk_L1_B233), .X(clk_L0_B3743));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R1_INV_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R2_INV_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R2_INV_1 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y34__R3_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3779));
  sky130_fd_sc_hd__clkbuf_4 T35Y35__R0_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3815));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R0_INV_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y35__R1_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3851));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R1_INV_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R2_INV_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R2_INV_1 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y35__R3_BUF_0 (.A(clk_L1_B242), .X(clk_L0_B3887));
  sky130_fd_sc_hd__clkbuf_4 T35Y36__R0_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3923));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R0_INV_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y36__R1_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3959));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R1_INV_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R2_INV_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R2_INV_1 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y36__R3_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3995));
  sky130_fd_sc_hd__clkbuf_4 T35Y37__R0_BUF_0 (.A(clk_L1_B251), .X(clk_L0_B4031));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R0_INV_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y37__R1_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4067));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R1_INV_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R2_INV_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R2_INV_1 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y37__R3_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4103));
  sky130_fd_sc_hd__clkbuf_4 T35Y38__R0_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4139));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R0_INV_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y38__R1_BUF_0 (.A(clk_L1_B260), .X(clk_L0_B4175));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R1_INV_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R2_INV_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R2_INV_1 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y38__R3_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4211));
  sky130_fd_sc_hd__clkbuf_4 T35Y39__R0_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4247));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R0_INV_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y39__R1_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4283));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R1_INV_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R2_INV_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R2_INV_1 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y39__R3_BUF_0 (.A(clk_L1_B269), .X(clk_L0_B4319));
  sky130_fd_sc_hd__clkbuf_4 T35Y3__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B9));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R0_INV_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y3__R1_BUF_0 (.A(clk_L1_B24), .X(clk_L0_B396));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R1_INV_0 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R2_INV_0 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R2_INV_1 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y3__R3_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B27));
  sky130_fd_sc_hd__clkbuf_4 T35Y40__R0_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4355));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R0_INV_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y40__R1_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4391));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R1_INV_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R2_INV_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R2_INV_1 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y40__R3_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4427));
  sky130_fd_sc_hd__clkbuf_4 T35Y41__R0_BUF_0 (.A(clk_L1_B278), .X(clk_L0_B4463));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R0_INV_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y41__R1_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4499));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R1_INV_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R2_INV_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R2_INV_1 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y41__R3_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4535));
  sky130_fd_sc_hd__clkbuf_4 T35Y42__R0_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4571));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R0_INV_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y42__R1_BUF_0 (.A(clk_L1_B287), .X(clk_L0_B4607));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R1_INV_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R2_INV_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R2_INV_1 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y42__R3_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4643));
  sky130_fd_sc_hd__clkbuf_4 T35Y43__R0_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4679));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R0_INV_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y43__R1_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4715));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R1_INV_0 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R2_INV_0 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R2_INV_1 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y43__R3_BUF_0 (.A(clk_L1_B296), .X(clk_L0_B4751));
  sky130_fd_sc_hd__clkbuf_4 T35Y44__R0_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4787));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R0_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y44__R1_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4823));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R1_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R2_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R2_INV_1 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y44__R3_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4859));
  sky130_fd_sc_hd__clkbuf_4 T35Y45__R0_BUF_0 (.A(clk_L1_B305), .X(clk_L0_B4895));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R0_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y45__R1_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4931));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R1_INV_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R2_INV_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R2_INV_1 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y45__R3_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4967));
  sky130_fd_sc_hd__clkbuf_4 T35Y46__R0_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5003));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R0_INV_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y46__R1_BUF_0 (.A(clk_L1_B314), .X(clk_L0_B5039));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R1_INV_0 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R2_INV_0 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R2_INV_1 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y46__R3_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5075));
  sky130_fd_sc_hd__clkbuf_4 T35Y47__R0_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5111));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R0_INV_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y47__R1_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5147));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R1_INV_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R2_INV_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R2_INV_1 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y47__R3_BUF_0 (.A(clk_L1_B323), .X(clk_L0_B5183));
  sky130_fd_sc_hd__clkbuf_4 T35Y48__R0_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5219));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R0_INV_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y48__R1_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5255));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R1_INV_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R2_INV_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R2_INV_1 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y48__R3_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5291));
  sky130_fd_sc_hd__clkbuf_4 T35Y49__R0_BUF_0 (.A(clk_L1_B332), .X(clk_L0_B5327));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R0_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y49__R1_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5363));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R1_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R2_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R2_INV_1 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y49__R3_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5399));
  sky130_fd_sc_hd__clkbuf_4 T35Y4__R0_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B468));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R0_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y4__R1_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B504));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R1_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R2_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R2_INV_1 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y4__R3_BUF_0 (.A(clk_L1_B33), .X(clk_L0_B540));
  sky130_fd_sc_hd__clkbuf_4 T35Y50__R0_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5435));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R0_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y50__R1_BUF_0 (.A(clk_L1_B341), .X(clk_L0_B5471));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R1_INV_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R2_INV_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R2_INV_1 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y50__R3_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5507));
  sky130_fd_sc_hd__clkbuf_4 T35Y51__R0_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5543));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R0_INV_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y51__R1_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5579));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R1_INV_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R2_INV_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R2_INV_1 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y51__R3_BUF_0 (.A(clk_L1_B350), .X(clk_L0_B5615));
  sky130_fd_sc_hd__clkbuf_4 T35Y52__R0_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5651));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R0_INV_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y52__R1_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5687));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R1_INV_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R2_INV_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R2_INV_1 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y52__R3_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5723));
  sky130_fd_sc_hd__clkbuf_4 T35Y53__R0_BUF_0 (.A(clk_L1_B359), .X(clk_L0_B5759));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R0_INV_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y53__R1_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5795));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R1_INV_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R2_INV_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R2_INV_1 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y53__R3_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5831));
  sky130_fd_sc_hd__clkbuf_4 T35Y54__R0_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5867));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R0_INV_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y54__R1_BUF_0 (.A(clk_L1_B368), .X(clk_L0_B5903));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R1_INV_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R2_INV_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R2_INV_1 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y54__R3_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5939));
  sky130_fd_sc_hd__clkbuf_4 T35Y55__R0_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5975));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R0_INV_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y55__R1_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6011));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R1_INV_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R2_INV_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R2_INV_1 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y55__R3_BUF_0 (.A(clk_L1_B377), .X(clk_L0_B6047));
  sky130_fd_sc_hd__clkbuf_4 T35Y56__R0_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6083));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R0_INV_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y56__R1_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6119));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R1_INV_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R2_INV_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R2_INV_1 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y56__R3_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6155));
  sky130_fd_sc_hd__clkbuf_4 T35Y57__R0_BUF_0 (.A(clk_L1_B386), .X(clk_L0_B6191));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R0_INV_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y57__R1_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6227));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R1_INV_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R2_INV_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R2_INV_1 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y57__R3_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6263));
  sky130_fd_sc_hd__clkbuf_4 T35Y58__R0_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6299));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R0_INV_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y58__R1_BUF_0 (.A(clk_L1_B395), .X(clk_L0_B6335));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R1_INV_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R2_INV_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R2_INV_1 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y58__R3_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6371));
  sky130_fd_sc_hd__clkbuf_4 T35Y59__R0_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6407));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R0_INV_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y59__R1_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6443));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R1_INV_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R2_INV_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R2_INV_1 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y59__R3_BUF_0 (.A(clk_L1_B404), .X(clk_L0_B6479));
  sky130_fd_sc_hd__clkbuf_4 T35Y5__R0_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B36));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R0_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y5__R1_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B612));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R1_INV_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R2_INV_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R2_INV_1 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y5__R3_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B648));
  sky130_fd_sc_hd__clkbuf_4 T35Y60__R0_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6515));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R0_INV_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y60__R1_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6551));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R1_INV_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R2_INV_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R2_INV_1 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y60__R3_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6587));
  sky130_fd_sc_hd__clkbuf_4 T35Y61__R0_BUF_0 (.A(clk_L1_B413), .X(clk_L0_B6623));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R0_INV_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y61__R1_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6659));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R1_INV_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R2_INV_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R2_INV_1 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y61__R3_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6695));
  sky130_fd_sc_hd__clkbuf_4 T35Y62__R0_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6731));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R0_INV_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y62__R1_BUF_0 (.A(clk_L1_B422), .X(clk_L0_B6767));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R1_INV_0 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R2_INV_0 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R2_INV_1 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y62__R3_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6803));
  sky130_fd_sc_hd__clkbuf_4 T35Y63__R0_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6839));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R0_INV_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y63__R1_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6875));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R1_INV_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R2_INV_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R2_INV_1 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y63__R3_BUF_0 (.A(clk_L1_B431), .X(clk_L0_B6911));
  sky130_fd_sc_hd__clkbuf_4 T35Y64__R0_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6947));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R0_INV_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y64__R1_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6983));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R1_INV_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R2_INV_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R2_INV_1 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y64__R3_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7019));
  sky130_fd_sc_hd__clkbuf_4 T35Y65__R0_BUF_0 (.A(clk_L1_B440), .X(clk_L0_B7055));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R0_INV_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y65__R1_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7091));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R1_INV_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R2_INV_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R2_INV_1 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y65__R3_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7127));
  sky130_fd_sc_hd__clkbuf_4 T35Y66__R0_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7163));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R0_INV_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y66__R1_BUF_0 (.A(clk_L1_B449), .X(clk_L0_B7199));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R1_INV_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R2_INV_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R2_INV_1 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y66__R3_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7235));
  sky130_fd_sc_hd__clkbuf_4 T35Y67__R0_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7271));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R0_INV_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y67__R1_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7307));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R1_INV_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R2_INV_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R2_INV_1 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y67__R3_BUF_0 (.A(clk_L1_B458), .X(clk_L0_B7343));
  sky130_fd_sc_hd__clkbuf_4 T35Y68__R0_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7379));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R0_INV_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y68__R1_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7415));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R1_INV_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R2_INV_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R2_INV_1 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y68__R3_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7451));
  sky130_fd_sc_hd__clkbuf_4 T35Y69__R0_BUF_0 (.A(clk_L1_B467), .X(clk_L0_B7487));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R0_INV_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y69__R1_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7523));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R1_INV_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R2_INV_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R2_INV_1 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y69__R3_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7559));
  sky130_fd_sc_hd__clkbuf_4 T35Y6__R0_BUF_0 (.A(clk_L1_B42), .X(clk_L0_B684));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R0_INV_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y6__R1_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B45));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R1_INV_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R2_INV_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R2_INV_1 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y6__R3_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B756));
  sky130_fd_sc_hd__clkbuf_4 T35Y70__R0_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7595));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R0_INV_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y70__R1_BUF_0 (.A(clk_L1_B476), .X(clk_L0_B7631));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R1_INV_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R2_INV_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R2_INV_1 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y70__R3_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7667));
  sky130_fd_sc_hd__clkbuf_4 T35Y71__R0_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7703));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R0_INV_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y71__R1_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7739));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R1_INV_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R2_INV_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R2_INV_1 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y71__R3_BUF_0 (.A(clk_L1_B485), .X(clk_L0_B7775));
  sky130_fd_sc_hd__clkbuf_4 T35Y72__R0_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7811));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R0_INV_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y72__R1_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7847));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R1_INV_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R2_INV_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R2_INV_1 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y72__R3_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7883));
  sky130_fd_sc_hd__clkbuf_4 T35Y73__R0_BUF_0 (.A(clk_L1_B494), .X(clk_L0_B7919));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R0_INV_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y73__R1_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7955));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R1_INV_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R2_INV_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R2_INV_1 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y73__R3_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7991));
  sky130_fd_sc_hd__clkbuf_4 T35Y74__R0_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8027));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R0_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y74__R1_BUF_0 (.A(clk_L1_B503), .X(clk_L0_B8063));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R1_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R2_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R2_INV_1 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y74__R3_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8099));
  sky130_fd_sc_hd__clkbuf_4 T35Y75__R0_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8135));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R0_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y75__R1_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8171));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R1_INV_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R2_INV_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R2_INV_1 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y75__R3_BUF_0 (.A(clk_L1_B512), .X(clk_L0_B8207));
  sky130_fd_sc_hd__clkbuf_4 T35Y76__R0_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8243));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R0_INV_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y76__R1_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8279));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R1_INV_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R2_INV_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R2_INV_1 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y76__R3_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8315));
  sky130_fd_sc_hd__clkbuf_4 T35Y77__R0_BUF_0 (.A(clk_L1_B521), .X(clk_L0_B8351));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R0_INV_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y77__R1_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8387));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R1_INV_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R2_INV_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R2_INV_1 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y77__R3_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8423));
  sky130_fd_sc_hd__clkbuf_4 T35Y78__R0_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8459));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R0_INV_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y78__R1_BUF_0 (.A(clk_L1_B530), .X(clk_L0_B8495));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R1_INV_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R2_INV_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R2_INV_1 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y78__R3_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8531));
  sky130_fd_sc_hd__clkbuf_4 T35Y79__R0_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8567));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R0_INV_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y79__R1_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8603));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R1_INV_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R2_INV_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R2_INV_1 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y79__R3_BUF_0 (.A(clk_L1_B539), .X(clk_L0_B8639));
  sky130_fd_sc_hd__clkbuf_4 T35Y7__R0_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B792));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R0_INV_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y7__R1_BUF_0 (.A(clk_L1_B51), .X(clk_L0_B828));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R1_INV_0 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R2_INV_0 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R2_INV_1 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y7__R3_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B54));
  sky130_fd_sc_hd__clkbuf_4 T35Y80__R0_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8675));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R0_INV_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y80__R1_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8711));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R1_INV_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R2_INV_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R2_INV_1 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y80__R3_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8747));
  sky130_fd_sc_hd__clkbuf_4 T35Y81__R0_BUF_0 (.A(clk_L1_B548), .X(clk_L0_B8783));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R0_INV_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y81__R1_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8819));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R1_INV_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R2_INV_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R2_INV_1 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y81__R3_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8855));
  sky130_fd_sc_hd__clkbuf_4 T35Y82__R0_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8891));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R0_INV_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y82__R1_BUF_0 (.A(clk_L1_B557), .X(clk_L0_B8927));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R1_INV_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R2_INV_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R2_INV_1 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y82__R3_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8963));
  sky130_fd_sc_hd__clkbuf_4 T35Y83__R0_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B8999));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R0_INV_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y83__R1_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9035));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R1_INV_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R2_INV_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R2_INV_1 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y83__R3_BUF_0 (.A(clk_L1_B566), .X(clk_L0_B9071));
  sky130_fd_sc_hd__clkbuf_4 T35Y84__R0_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9107));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R0_INV_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y84__R1_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9143));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R1_INV_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R2_INV_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R2_INV_1 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y84__R3_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9179));
  sky130_fd_sc_hd__clkbuf_4 T35Y85__R0_BUF_0 (.A(clk_L1_B575), .X(clk_L0_B9215));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R0_INV_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y85__R1_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9251));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R1_INV_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R2_INV_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R2_INV_1 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y85__R3_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9287));
  sky130_fd_sc_hd__clkbuf_4 T35Y86__R0_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9323));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R0_INV_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y86__R1_BUF_0 (.A(clk_L1_B584), .X(clk_L0_B9359));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R1_INV_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R2_INV_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R2_INV_1 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y86__R3_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9395));
  sky130_fd_sc_hd__clkbuf_4 T35Y87__R0_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9431));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R0_INV_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y87__R1_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9467));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R1_INV_0 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R2_INV_0 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R2_INV_1 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y87__R3_BUF_0 (.A(clk_L1_B593), .X(clk_L0_B9503));
  sky130_fd_sc_hd__clkbuf_4 T35Y88__R0_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9539));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R0_INV_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y88__R1_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9575));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R1_INV_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R2_INV_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R2_INV_1 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y88__R3_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9611));
  sky130_fd_sc_hd__clkbuf_4 T35Y89__R0_BUF_0 (.A(clk_L1_B602), .X(clk_L0_B9647));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R0_INV_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y89__R1_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9683));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R1_INV_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R2_INV_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R2_INV_1 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y89__R3_BUF_0 (.A(clk_L1_B607), .X(clk_L0_B9719));
  sky130_fd_sc_hd__clkbuf_4 T35Y8__R0_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B900));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R0_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y8__R1_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B936));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R1_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R2_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R2_INV_1 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y8__R3_BUF_0 (.A(clk_L1_B60), .X(clk_L0_B972));
  sky130_fd_sc_hd__clkbuf_4 T35Y9__R0_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B63));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R0_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y9__R1_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1044));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R1_INV_0 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R2_INV_0 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R2_INV_1 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y9__R3_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1080));
  sky130_fd_sc_hd__clkbuf_4 T3Y0__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B13));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R0_INV_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y0__R1_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B3));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R1_INV_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R2_INV_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R2_INV_1 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B83));
  sky130_fd_sc_hd__clkbuf_4 T3Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1084));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R0_INV_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y10__R1_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B70));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R1_INV_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R2_INV_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R2_INV_1 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1156));
  sky130_fd_sc_hd__clkbuf_4 T3Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1192));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R0_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1228));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R1_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R2_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R2_INV_1 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y11__R3_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B79));
  sky130_fd_sc_hd__clkbuf_4 T3Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1300));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R0_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1336));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R1_INV_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R2_INV_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R2_INV_1 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1372));
  sky130_fd_sc_hd__clkbuf_4 T3Y13__R0_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B88));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R0_INV_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1444));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R1_INV_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R2_INV_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R2_INV_1 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1480));
  sky130_fd_sc_hd__clkbuf_4 T3Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1516));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R0_INV_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y14__R1_BUF_0 (.A(clk_L1_B96), .X(clk_L0_B1551));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R1_INV_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R2_INV_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R2_INV_1 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1587));
  sky130_fd_sc_hd__clkbuf_4 T3Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1623));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R0_INV_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1659));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R1_INV_0 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R2_INV_0 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R2_INV_1 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y15__R3_BUF_0 (.A(clk_L1_B105), .X(clk_L0_B1695));
  sky130_fd_sc_hd__clkbuf_4 T3Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1731));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R0_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1767));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R1_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R2_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R2_INV_1 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1803));
  sky130_fd_sc_hd__clkbuf_4 T3Y17__R0_BUF_0 (.A(clk_L1_B114), .X(clk_L0_B1839));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R0_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1875));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R1_INV_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R2_INV_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R2_INV_1 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1911));
  sky130_fd_sc_hd__clkbuf_4 T3Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1947));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R0_INV_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y18__R1_BUF_0 (.A(clk_L1_B123), .X(clk_L0_B1983));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R1_INV_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R2_INV_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R2_INV_1 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2019));
  sky130_fd_sc_hd__clkbuf_4 T3Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2055));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R0_INV_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2091));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R1_INV_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R2_INV_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R2_INV_1 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y19__R3_BUF_0 (.A(clk_L1_B132), .X(clk_L0_B2127));
  sky130_fd_sc_hd__clkbuf_4 T3Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B118));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R0_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B153));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R1_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R2_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R2_INV_1 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B188));
  sky130_fd_sc_hd__clkbuf_4 T3Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2163));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R0_INV_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2199));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R1_INV_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R2_INV_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R2_INV_1 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2235));
  sky130_fd_sc_hd__clkbuf_4 T3Y21__R0_BUF_0 (.A(clk_L1_B141), .X(clk_L0_B2271));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R0_INV_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2307));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R1_INV_0 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R2_INV_0 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R2_INV_1 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2343));
  sky130_fd_sc_hd__clkbuf_4 T3Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2379));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R0_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y22__R1_BUF_0 (.A(clk_L1_B150), .X(clk_L0_B2415));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R1_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R2_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R2_INV_1 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2451));
  sky130_fd_sc_hd__clkbuf_4 T3Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2487));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R0_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2523));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R1_INV_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R2_INV_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R2_INV_1 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y23__R3_BUF_0 (.A(clk_L1_B159), .X(clk_L0_B2559));
  sky130_fd_sc_hd__clkbuf_4 T3Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2595));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R0_INV_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2631));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R1_INV_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R2_INV_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R2_INV_1 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2667));
  sky130_fd_sc_hd__clkbuf_4 T3Y25__R0_BUF_0 (.A(clk_L1_B168), .X(clk_L0_B2703));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R0_INV_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2739));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R1_INV_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R2_INV_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R2_INV_1 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2775));
  sky130_fd_sc_hd__clkbuf_4 T3Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2811));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R0_INV_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y26__R1_BUF_0 (.A(clk_L1_B177), .X(clk_L0_B2847));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R1_INV_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R2_INV_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R2_INV_1 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2883));
  sky130_fd_sc_hd__clkbuf_4 T3Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2919));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R0_INV_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2955));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R1_INV_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R2_INV_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R2_INV_1 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y27__R3_BUF_0 (.A(clk_L1_B186), .X(clk_L0_B2991));
  sky130_fd_sc_hd__clkbuf_4 T3Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3027));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R0_INV_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3063));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R1_INV_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R2_INV_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R2_INV_1 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3099));
  sky130_fd_sc_hd__clkbuf_4 T3Y29__R0_BUF_0 (.A(clk_L1_B195), .X(clk_L0_B3135));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R0_INV_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3171));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R1_INV_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R2_INV_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R2_INV_1 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3207));
  sky130_fd_sc_hd__clkbuf_4 T3Y2__R0_BUF_0 (.A(clk_L1_B13), .X(clk_L0_B223));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R0_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B258));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R1_INV_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R2_INV_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R2_INV_1 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B294));
  sky130_fd_sc_hd__clkbuf_4 T3Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3243));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R0_INV_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y30__R1_BUF_0 (.A(clk_L1_B204), .X(clk_L0_B3279));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R1_INV_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R2_INV_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R2_INV_1 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3315));
  sky130_fd_sc_hd__clkbuf_4 T3Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3351));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R0_INV_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3387));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R1_INV_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R2_INV_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R2_INV_1 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y31__R3_BUF_0 (.A(clk_L1_B213), .X(clk_L0_B3423));
  sky130_fd_sc_hd__clkbuf_4 T3Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3459));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R0_INV_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3495));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R1_INV_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R2_INV_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R2_INV_1 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3531));
  sky130_fd_sc_hd__clkbuf_4 T3Y33__R0_BUF_0 (.A(clk_L1_B222), .X(clk_L0_B3567));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R0_INV_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3603));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R1_INV_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R2_INV_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R2_INV_1 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3639));
  sky130_fd_sc_hd__clkbuf_4 T3Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3675));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R0_INV_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y34__R1_BUF_0 (.A(clk_L1_B231), .X(clk_L0_B3711));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R1_INV_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R2_INV_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R2_INV_1 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3747));
  sky130_fd_sc_hd__clkbuf_4 T3Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3783));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R0_INV_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3819));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R1_INV_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R2_INV_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R2_INV_1 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y35__R3_BUF_0 (.A(clk_L1_B240), .X(clk_L0_B3855));
  sky130_fd_sc_hd__clkbuf_4 T3Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3891));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R0_INV_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3927));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R1_INV_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R2_INV_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R2_INV_1 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3963));
  sky130_fd_sc_hd__clkbuf_4 T3Y37__R0_BUF_0 (.A(clk_L1_B249), .X(clk_L0_B3999));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R0_INV_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4035));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R1_INV_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R2_INV_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R2_INV_1 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4071));
  sky130_fd_sc_hd__clkbuf_4 T3Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4107));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R0_INV_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y38__R1_BUF_0 (.A(clk_L1_B258), .X(clk_L0_B4143));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R1_INV_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R2_INV_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R2_INV_1 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4179));
  sky130_fd_sc_hd__clkbuf_4 T3Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4215));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R0_INV_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4251));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R1_INV_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R2_INV_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R2_INV_1 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y39__R3_BUF_0 (.A(clk_L1_B267), .X(clk_L0_B4287));
  sky130_fd_sc_hd__clkbuf_4 T3Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B329));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R0_INV_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B364));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R1_INV_0 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R2_INV_0 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R2_INV_1 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y3__R3_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B25));
  sky130_fd_sc_hd__clkbuf_4 T3Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4323));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R0_INV_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4359));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R1_INV_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R2_INV_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R2_INV_1 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4395));
  sky130_fd_sc_hd__clkbuf_4 T3Y41__R0_BUF_0 (.A(clk_L1_B276), .X(clk_L0_B4431));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R0_INV_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4467));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R1_INV_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R2_INV_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R2_INV_1 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4503));
  sky130_fd_sc_hd__clkbuf_4 T3Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4539));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R0_INV_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y42__R1_BUF_0 (.A(clk_L1_B285), .X(clk_L0_B4575));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R1_INV_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R2_INV_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R2_INV_1 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4611));
  sky130_fd_sc_hd__clkbuf_4 T3Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4647));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R0_INV_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4683));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R1_INV_0 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R2_INV_0 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R2_INV_1 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y43__R3_BUF_0 (.A(clk_L1_B294), .X(clk_L0_B4719));
  sky130_fd_sc_hd__clkbuf_4 T3Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4755));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R0_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4791));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R1_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R2_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R2_INV_1 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4827));
  sky130_fd_sc_hd__clkbuf_4 T3Y45__R0_BUF_0 (.A(clk_L1_B303), .X(clk_L0_B4863));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R0_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4899));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R1_INV_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R2_INV_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R2_INV_1 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4935));
  sky130_fd_sc_hd__clkbuf_4 T3Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4971));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R0_INV_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y46__R1_BUF_0 (.A(clk_L1_B312), .X(clk_L0_B5007));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R1_INV_0 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R2_INV_0 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R2_INV_1 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5043));
  sky130_fd_sc_hd__clkbuf_4 T3Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5079));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R0_INV_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5115));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R1_INV_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R2_INV_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R2_INV_1 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y47__R3_BUF_0 (.A(clk_L1_B321), .X(clk_L0_B5151));
  sky130_fd_sc_hd__clkbuf_4 T3Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5187));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R0_INV_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5223));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R1_INV_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R2_INV_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R2_INV_1 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5259));
  sky130_fd_sc_hd__clkbuf_4 T3Y49__R0_BUF_0 (.A(clk_L1_B330), .X(clk_L0_B5295));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R0_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5331));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R1_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R2_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R2_INV_1 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5367));
  sky130_fd_sc_hd__clkbuf_4 T3Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B436));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R0_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B472));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R1_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R2_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R2_INV_1 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B508));
  sky130_fd_sc_hd__clkbuf_4 T3Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5403));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R0_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y50__R1_BUF_0 (.A(clk_L1_B339), .X(clk_L0_B5439));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R1_INV_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R2_INV_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R2_INV_1 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5475));
  sky130_fd_sc_hd__clkbuf_4 T3Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5511));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R0_INV_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5547));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R1_INV_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R2_INV_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R2_INV_1 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y51__R3_BUF_0 (.A(clk_L1_B348), .X(clk_L0_B5583));
  sky130_fd_sc_hd__clkbuf_4 T3Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5619));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R0_INV_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5655));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R1_INV_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R2_INV_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R2_INV_1 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5691));
  sky130_fd_sc_hd__clkbuf_4 T3Y53__R0_BUF_0 (.A(clk_L1_B357), .X(clk_L0_B5727));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R0_INV_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5763));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R1_INV_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R2_INV_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R2_INV_1 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5799));
  sky130_fd_sc_hd__clkbuf_4 T3Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5835));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R0_INV_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y54__R1_BUF_0 (.A(clk_L1_B366), .X(clk_L0_B5871));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R1_INV_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R2_INV_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R2_INV_1 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5907));
  sky130_fd_sc_hd__clkbuf_4 T3Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5943));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R0_INV_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5979));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R1_INV_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R2_INV_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R2_INV_1 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y55__R3_BUF_0 (.A(clk_L1_B375), .X(clk_L0_B6015));
  sky130_fd_sc_hd__clkbuf_4 T3Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6051));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R0_INV_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6087));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R1_INV_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R2_INV_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R2_INV_1 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6123));
  sky130_fd_sc_hd__clkbuf_4 T3Y57__R0_BUF_0 (.A(clk_L1_B384), .X(clk_L0_B6159));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R0_INV_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6195));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R1_INV_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R2_INV_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R2_INV_1 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6231));
  sky130_fd_sc_hd__clkbuf_4 T3Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6267));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R0_INV_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y58__R1_BUF_0 (.A(clk_L1_B393), .X(clk_L0_B6303));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R1_INV_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R2_INV_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R2_INV_1 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6339));
  sky130_fd_sc_hd__clkbuf_4 T3Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6375));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R0_INV_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6411));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R1_INV_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R2_INV_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R2_INV_1 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y59__R3_BUF_0 (.A(clk_L1_B402), .X(clk_L0_B6447));
  sky130_fd_sc_hd__clkbuf_4 T3Y5__R0_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B34));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R0_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B580));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R1_INV_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R2_INV_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R2_INV_1 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B616));
  sky130_fd_sc_hd__clkbuf_4 T3Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6483));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R0_INV_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6519));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R1_INV_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R2_INV_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R2_INV_1 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6555));
  sky130_fd_sc_hd__clkbuf_4 T3Y61__R0_BUF_0 (.A(clk_L1_B411), .X(clk_L0_B6591));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R0_INV_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6627));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R1_INV_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R2_INV_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R2_INV_1 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6663));
  sky130_fd_sc_hd__clkbuf_4 T3Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6699));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R0_INV_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y62__R1_BUF_0 (.A(clk_L1_B420), .X(clk_L0_B6735));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R1_INV_0 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R2_INV_0 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R2_INV_1 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6771));
  sky130_fd_sc_hd__clkbuf_4 T3Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6807));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R0_INV_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6843));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R1_INV_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R2_INV_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R2_INV_1 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y63__R3_BUF_0 (.A(clk_L1_B429), .X(clk_L0_B6879));
  sky130_fd_sc_hd__clkbuf_4 T3Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6915));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R0_INV_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6951));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R1_INV_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R2_INV_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R2_INV_1 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6987));
  sky130_fd_sc_hd__clkbuf_4 T3Y65__R0_BUF_0 (.A(clk_L1_B438), .X(clk_L0_B7023));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R0_INV_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7059));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R1_INV_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R2_INV_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R2_INV_1 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7095));
  sky130_fd_sc_hd__clkbuf_4 T3Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7131));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R0_INV_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y66__R1_BUF_0 (.A(clk_L1_B447), .X(clk_L0_B7167));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R1_INV_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R2_INV_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R2_INV_1 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7203));
  sky130_fd_sc_hd__clkbuf_4 T3Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7239));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R0_INV_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7275));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R1_INV_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R2_INV_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R2_INV_1 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y67__R3_BUF_0 (.A(clk_L1_B456), .X(clk_L0_B7311));
  sky130_fd_sc_hd__clkbuf_4 T3Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7347));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R0_INV_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7383));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R1_INV_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R2_INV_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R2_INV_1 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7419));
  sky130_fd_sc_hd__clkbuf_4 T3Y69__R0_BUF_0 (.A(clk_L1_B465), .X(clk_L0_B7455));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R0_INV_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7491));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R1_INV_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R2_INV_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R2_INV_1 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7527));
  sky130_fd_sc_hd__clkbuf_4 T3Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B652));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R0_INV_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y6__R1_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B43));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R1_INV_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R2_INV_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R2_INV_1 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B724));
  sky130_fd_sc_hd__clkbuf_4 T3Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7563));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R0_INV_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y70__R1_BUF_0 (.A(clk_L1_B474), .X(clk_L0_B7599));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R1_INV_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R2_INV_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R2_INV_1 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7635));
  sky130_fd_sc_hd__clkbuf_4 T3Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7671));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R0_INV_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7707));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R1_INV_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R2_INV_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R2_INV_1 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y71__R3_BUF_0 (.A(clk_L1_B483), .X(clk_L0_B7743));
  sky130_fd_sc_hd__clkbuf_4 T3Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7779));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R0_INV_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7815));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R1_INV_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R2_INV_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R2_INV_1 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7851));
  sky130_fd_sc_hd__clkbuf_4 T3Y73__R0_BUF_0 (.A(clk_L1_B492), .X(clk_L0_B7887));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R0_INV_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7923));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R1_INV_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R2_INV_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R2_INV_1 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7959));
  sky130_fd_sc_hd__clkbuf_4 T3Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7995));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R0_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y74__R1_BUF_0 (.A(clk_L1_B501), .X(clk_L0_B8031));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R1_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R2_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R2_INV_1 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8067));
  sky130_fd_sc_hd__clkbuf_4 T3Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8103));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R0_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8139));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R1_INV_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R2_INV_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R2_INV_1 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y75__R3_BUF_0 (.A(clk_L1_B510), .X(clk_L0_B8175));
  sky130_fd_sc_hd__clkbuf_4 T3Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8211));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R0_INV_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8247));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R1_INV_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R2_INV_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R2_INV_1 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8283));
  sky130_fd_sc_hd__clkbuf_4 T3Y77__R0_BUF_0 (.A(clk_L1_B519), .X(clk_L0_B8319));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R0_INV_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8355));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R1_INV_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R2_INV_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R2_INV_1 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8391));
  sky130_fd_sc_hd__clkbuf_4 T3Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8427));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R0_INV_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y78__R1_BUF_0 (.A(clk_L1_B528), .X(clk_L0_B8463));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R1_INV_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R2_INV_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R2_INV_1 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8499));
  sky130_fd_sc_hd__clkbuf_4 T3Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8535));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R0_INV_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8571));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R1_INV_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R2_INV_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R2_INV_1 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y79__R3_BUF_0 (.A(clk_L1_B537), .X(clk_L0_B8607));
  sky130_fd_sc_hd__clkbuf_4 T3Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B760));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R0_INV_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B796));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R1_INV_0 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R2_INV_0 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R2_INV_1 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y7__R3_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B52));
  sky130_fd_sc_hd__clkbuf_4 T3Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8643));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R0_INV_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8679));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R1_INV_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R2_INV_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R2_INV_1 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8715));
  sky130_fd_sc_hd__clkbuf_4 T3Y81__R0_BUF_0 (.A(clk_L1_B546), .X(clk_L0_B8751));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R0_INV_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8787));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R1_INV_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R2_INV_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R2_INV_1 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8823));
  sky130_fd_sc_hd__clkbuf_4 T3Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8859));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R0_INV_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y82__R1_BUF_0 (.A(clk_L1_B555), .X(clk_L0_B8895));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R1_INV_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R2_INV_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R2_INV_1 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8931));
  sky130_fd_sc_hd__clkbuf_4 T3Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8967));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R0_INV_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9003));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R1_INV_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R2_INV_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R2_INV_1 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y83__R3_BUF_0 (.A(clk_L1_B564), .X(clk_L0_B9039));
  sky130_fd_sc_hd__clkbuf_4 T3Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9075));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R0_INV_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9111));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R1_INV_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R2_INV_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R2_INV_1 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9147));
  sky130_fd_sc_hd__clkbuf_4 T3Y85__R0_BUF_0 (.A(clk_L1_B573), .X(clk_L0_B9183));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R0_INV_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9219));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R1_INV_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R2_INV_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R2_INV_1 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9255));
  sky130_fd_sc_hd__clkbuf_4 T3Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9291));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R0_INV_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y86__R1_BUF_0 (.A(clk_L1_B582), .X(clk_L0_B9327));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R1_INV_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R2_INV_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R2_INV_1 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9363));
  sky130_fd_sc_hd__clkbuf_4 T3Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9399));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R0_INV_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9435));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R1_INV_0 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R2_INV_0 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R2_INV_1 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y87__R3_BUF_0 (.A(clk_L1_B591), .X(clk_L0_B9471));
  sky130_fd_sc_hd__clkbuf_4 T3Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9507));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R0_INV_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9543));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R1_INV_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R2_INV_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R2_INV_1 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9579));
  sky130_fd_sc_hd__clkbuf_4 T3Y89__R0_BUF_0 (.A(clk_L1_B600), .X(clk_L0_B9615));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R0_INV_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9651));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R1_INV_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R2_INV_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R2_INV_1 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9687));
  sky130_fd_sc_hd__clkbuf_4 T3Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B868));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R0_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B904));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R1_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R2_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R2_INV_1 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B940));
  sky130_fd_sc_hd__clkbuf_4 T3Y9__R0_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B61));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R0_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1012));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R1_INV_0 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R2_INV_0 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R2_INV_1 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1048));
  sky130_fd_sc_hd__clkbuf_4 T4Y0__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B14));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R0_INV_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B49));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R1_INV_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R2_INV_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R2_INV_1 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B84));
  sky130_fd_sc_hd__clkbuf_4 T4Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1085));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R0_INV_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1121));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R1_INV_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R2_INV_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R2_INV_1 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1157));
  sky130_fd_sc_hd__clkbuf_4 T4Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1193));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R0_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1229));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R1_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R2_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R2_INV_1 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1265));
  sky130_fd_sc_hd__clkbuf_4 T4Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1301));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R0_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1337));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R1_INV_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R2_INV_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R2_INV_1 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1373));
  sky130_fd_sc_hd__clkbuf_4 T4Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1409));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R0_INV_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1445));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R1_INV_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R2_INV_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R2_INV_1 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1481));
  sky130_fd_sc_hd__clkbuf_4 T4Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1517));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R0_INV_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y14__R1_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B97));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R1_INV_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R2_INV_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R2_INV_1 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1588));
  sky130_fd_sc_hd__clkbuf_4 T4Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1624));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R0_INV_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1660));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R1_INV_0 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R2_INV_0 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R2_INV_1 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y15__R3_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B106));
  sky130_fd_sc_hd__clkbuf_4 T4Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1732));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R0_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1768));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R1_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R2_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R2_INV_1 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1804));
  sky130_fd_sc_hd__clkbuf_4 T4Y17__R0_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B115));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R0_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1876));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R1_INV_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R2_INV_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R2_INV_1 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1912));
  sky130_fd_sc_hd__clkbuf_4 T4Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1948));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R0_INV_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y18__R1_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B124));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R1_INV_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R2_INV_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R2_INV_1 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2020));
  sky130_fd_sc_hd__clkbuf_4 T4Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2056));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R0_INV_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2092));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R1_INV_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R2_INV_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R2_INV_1 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y19__R3_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B133));
  sky130_fd_sc_hd__clkbuf_4 T4Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B119));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R0_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B154));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R1_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R2_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R2_INV_1 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B189));
  sky130_fd_sc_hd__clkbuf_4 T4Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2164));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R0_INV_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2200));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R1_INV_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R2_INV_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R2_INV_1 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2236));
  sky130_fd_sc_hd__clkbuf_4 T4Y21__R0_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B142));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R0_INV_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2308));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R1_INV_0 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R2_INV_0 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R2_INV_1 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2344));
  sky130_fd_sc_hd__clkbuf_4 T4Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2380));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R0_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y22__R1_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B151));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R1_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R2_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R2_INV_1 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2452));
  sky130_fd_sc_hd__clkbuf_4 T4Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2488));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R0_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2524));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R1_INV_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R2_INV_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R2_INV_1 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y23__R3_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B10));
  sky130_fd_sc_hd__clkbuf_4 T4Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2596));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R0_INV_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2632));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R1_INV_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R2_INV_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R2_INV_1 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2668));
  sky130_fd_sc_hd__clkbuf_4 T4Y25__R0_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B169));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R0_INV_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2740));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R1_INV_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R2_INV_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R2_INV_1 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2776));
  sky130_fd_sc_hd__clkbuf_4 T4Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2812));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R0_INV_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y26__R1_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B178));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R1_INV_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R2_INV_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R2_INV_1 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2884));
  sky130_fd_sc_hd__clkbuf_4 T4Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2920));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R0_INV_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2956));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R1_INV_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R2_INV_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R2_INV_1 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y27__R3_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B187));
  sky130_fd_sc_hd__clkbuf_4 T4Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3028));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R0_INV_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3064));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R1_INV_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R2_INV_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R2_INV_1 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3100));
  sky130_fd_sc_hd__clkbuf_4 T4Y29__R0_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B196));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R0_INV_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3172));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R1_INV_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R2_INV_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R2_INV_1 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3208));
  sky130_fd_sc_hd__clkbuf_4 T4Y2__R0_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B14));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R0_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B259));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R1_INV_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R2_INV_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R2_INV_1 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B295));
  sky130_fd_sc_hd__clkbuf_4 T4Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3244));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R0_INV_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y30__R1_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B205));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R1_INV_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R2_INV_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R2_INV_1 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3316));
  sky130_fd_sc_hd__clkbuf_4 T4Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3352));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R0_INV_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3388));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R1_INV_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R2_INV_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R2_INV_1 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y31__R3_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B214));
  sky130_fd_sc_hd__clkbuf_4 T4Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3460));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R0_INV_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3496));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R1_INV_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R2_INV_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R2_INV_1 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3532));
  sky130_fd_sc_hd__clkbuf_4 T4Y33__R0_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B223));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R0_INV_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3604));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R1_INV_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R2_INV_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R2_INV_1 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3640));
  sky130_fd_sc_hd__clkbuf_4 T4Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3676));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R0_INV_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y34__R1_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B232));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R1_INV_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R2_INV_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R2_INV_1 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3748));
  sky130_fd_sc_hd__clkbuf_4 T4Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3784));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R0_INV_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3820));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R1_INV_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R2_INV_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R2_INV_1 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y35__R3_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B241));
  sky130_fd_sc_hd__clkbuf_4 T4Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3892));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R0_INV_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3928));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R1_INV_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R2_INV_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R2_INV_1 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3964));
  sky130_fd_sc_hd__clkbuf_4 T4Y37__R0_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B250));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R0_INV_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4036));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R1_INV_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R2_INV_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R2_INV_1 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4072));
  sky130_fd_sc_hd__clkbuf_4 T4Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4108));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R0_INV_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y38__R1_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B259));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R1_INV_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R2_INV_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R2_INV_1 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4180));
  sky130_fd_sc_hd__clkbuf_4 T4Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4216));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R0_INV_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4252));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R1_INV_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R2_INV_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R2_INV_1 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y39__R3_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B268));
  sky130_fd_sc_hd__clkbuf_4 T4Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B330));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R0_INV_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B365));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R1_INV_0 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R2_INV_0 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R2_INV_1 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B401));
  sky130_fd_sc_hd__clkbuf_4 T4Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4324));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R0_INV_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4360));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R1_INV_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R2_INV_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R2_INV_1 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4396));
  sky130_fd_sc_hd__clkbuf_4 T4Y41__R0_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B277));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R0_INV_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4468));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R1_INV_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R2_INV_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R2_INV_1 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4504));
  sky130_fd_sc_hd__clkbuf_4 T4Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4540));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R0_INV_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y42__R1_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B286));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R1_INV_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R2_INV_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R2_INV_1 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4612));
  sky130_fd_sc_hd__clkbuf_4 T4Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4648));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R0_INV_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4684));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R1_INV_0 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R2_INV_0 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R2_INV_1 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y43__R3_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B295));
  sky130_fd_sc_hd__clkbuf_4 T4Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4756));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R0_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4792));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R1_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R2_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R2_INV_1 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4828));
  sky130_fd_sc_hd__clkbuf_4 T4Y45__R0_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B19));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R0_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4900));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R1_INV_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R2_INV_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R2_INV_1 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4936));
  sky130_fd_sc_hd__clkbuf_4 T4Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4972));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R0_INV_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y46__R1_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B313));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R1_INV_0 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R2_INV_0 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R2_INV_1 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5044));
  sky130_fd_sc_hd__clkbuf_4 T4Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5080));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R0_INV_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5116));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R1_INV_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R2_INV_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R2_INV_1 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y47__R3_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B322));
  sky130_fd_sc_hd__clkbuf_4 T4Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5188));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R0_INV_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5224));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R1_INV_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R2_INV_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R2_INV_1 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5260));
  sky130_fd_sc_hd__clkbuf_4 T4Y49__R0_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B331));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R0_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5332));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R1_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R2_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R2_INV_1 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5368));
  sky130_fd_sc_hd__clkbuf_4 T4Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B437));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R0_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B473));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R1_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R2_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R2_INV_1 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B509));
  sky130_fd_sc_hd__clkbuf_4 T4Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5404));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R0_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y50__R1_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B340));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R1_INV_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R2_INV_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R2_INV_1 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5476));
  sky130_fd_sc_hd__clkbuf_4 T4Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5512));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R0_INV_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5548));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R1_INV_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R2_INV_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R2_INV_1 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y51__R3_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B349));
  sky130_fd_sc_hd__clkbuf_4 T4Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5620));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R0_INV_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5656));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R1_INV_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R2_INV_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R2_INV_1 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5692));
  sky130_fd_sc_hd__clkbuf_4 T4Y53__R0_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B358));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R0_INV_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5764));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R1_INV_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R2_INV_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R2_INV_1 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5800));
  sky130_fd_sc_hd__clkbuf_4 T4Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5836));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R0_INV_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y54__R1_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B367));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R1_INV_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R2_INV_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R2_INV_1 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5908));
  sky130_fd_sc_hd__clkbuf_4 T4Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5944));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R0_INV_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5980));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R1_INV_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R2_INV_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R2_INV_1 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y55__R3_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B376));
  sky130_fd_sc_hd__clkbuf_4 T4Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6052));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R0_INV_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6088));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R1_INV_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R2_INV_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R2_INV_1 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6124));
  sky130_fd_sc_hd__clkbuf_4 T4Y57__R0_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B385));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R0_INV_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6196));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R1_INV_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R2_INV_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R2_INV_1 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6232));
  sky130_fd_sc_hd__clkbuf_4 T4Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6268));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R0_INV_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y58__R1_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B394));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R1_INV_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R2_INV_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R2_INV_1 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6340));
  sky130_fd_sc_hd__clkbuf_4 T4Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6376));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R0_INV_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6412));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R1_INV_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R2_INV_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R2_INV_1 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y59__R3_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B403));
  sky130_fd_sc_hd__clkbuf_4 T4Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B545));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R0_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B581));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R1_INV_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R2_INV_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R2_INV_1 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B617));
  sky130_fd_sc_hd__clkbuf_4 T4Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6484));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R0_INV_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6520));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R1_INV_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R2_INV_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R2_INV_1 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6556));
  sky130_fd_sc_hd__clkbuf_4 T4Y61__R0_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B412));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R0_INV_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6628));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R1_INV_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R2_INV_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R2_INV_1 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6664));
  sky130_fd_sc_hd__clkbuf_4 T4Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6700));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R0_INV_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y62__R1_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B421));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R1_INV_0 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R2_INV_0 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R2_INV_1 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6772));
  sky130_fd_sc_hd__clkbuf_4 T4Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6808));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R0_INV_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6844));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R1_INV_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R2_INV_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R2_INV_1 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y63__R3_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B430));
  sky130_fd_sc_hd__clkbuf_4 T4Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6916));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R0_INV_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6952));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R1_INV_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R2_INV_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R2_INV_1 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6988));
  sky130_fd_sc_hd__clkbuf_4 T4Y65__R0_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B439));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R0_INV_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7060));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R1_INV_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R2_INV_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R2_INV_1 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7096));
  sky130_fd_sc_hd__clkbuf_4 T4Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7132));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R0_INV_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y66__R1_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B28));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R1_INV_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R2_INV_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R2_INV_1 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7204));
  sky130_fd_sc_hd__clkbuf_4 T4Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7240));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R0_INV_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7276));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R1_INV_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R2_INV_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R2_INV_1 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y67__R3_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B457));
  sky130_fd_sc_hd__clkbuf_4 T4Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7348));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R0_INV_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7384));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R1_INV_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R2_INV_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R2_INV_1 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7420));
  sky130_fd_sc_hd__clkbuf_4 T4Y69__R0_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B466));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R0_INV_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7492));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R1_INV_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R2_INV_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R2_INV_1 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7528));
  sky130_fd_sc_hd__clkbuf_4 T4Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B653));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R0_INV_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B689));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R1_INV_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R2_INV_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R2_INV_1 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B725));
  sky130_fd_sc_hd__clkbuf_4 T4Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7564));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R0_INV_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y70__R1_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B475));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R1_INV_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R2_INV_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R2_INV_1 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7636));
  sky130_fd_sc_hd__clkbuf_4 T4Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7672));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R0_INV_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7708));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R1_INV_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R2_INV_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R2_INV_1 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y71__R3_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B484));
  sky130_fd_sc_hd__clkbuf_4 T4Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7780));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R0_INV_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7816));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R1_INV_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R2_INV_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R2_INV_1 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7852));
  sky130_fd_sc_hd__clkbuf_4 T4Y73__R0_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B493));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R0_INV_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7924));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R1_INV_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R2_INV_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R2_INV_1 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7960));
  sky130_fd_sc_hd__clkbuf_4 T4Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7996));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R0_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y74__R1_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B502));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R1_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R2_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R2_INV_1 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8068));
  sky130_fd_sc_hd__clkbuf_4 T4Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8104));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R0_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8140));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R1_INV_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R2_INV_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R2_INV_1 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y75__R3_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B511));
  sky130_fd_sc_hd__clkbuf_4 T4Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8212));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R0_INV_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8248));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R1_INV_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R2_INV_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R2_INV_1 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8284));
  sky130_fd_sc_hd__clkbuf_4 T4Y77__R0_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B520));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R0_INV_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8356));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R1_INV_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R2_INV_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R2_INV_1 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8392));
  sky130_fd_sc_hd__clkbuf_4 T4Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8428));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R0_INV_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y78__R1_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B529));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R1_INV_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R2_INV_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R2_INV_1 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8500));
  sky130_fd_sc_hd__clkbuf_4 T4Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8536));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R0_INV_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8572));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R1_INV_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R2_INV_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R2_INV_1 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y79__R3_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B538));
  sky130_fd_sc_hd__clkbuf_4 T4Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B761));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R0_INV_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B797));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R1_INV_0 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R2_INV_0 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R2_INV_1 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B833));
  sky130_fd_sc_hd__clkbuf_4 T4Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8644));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R0_INV_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8680));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R1_INV_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R2_INV_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R2_INV_1 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8716));
  sky130_fd_sc_hd__clkbuf_4 T4Y81__R0_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B547));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R0_INV_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8788));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R1_INV_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R2_INV_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R2_INV_1 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8824));
  sky130_fd_sc_hd__clkbuf_4 T4Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8860));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R0_INV_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y82__R1_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B556));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R1_INV_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R2_INV_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R2_INV_1 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8932));
  sky130_fd_sc_hd__clkbuf_4 T4Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8968));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R0_INV_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9004));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R1_INV_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R2_INV_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R2_INV_1 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y83__R3_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B565));
  sky130_fd_sc_hd__clkbuf_4 T4Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9076));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R0_INV_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9112));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R1_INV_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R2_INV_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R2_INV_1 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9148));
  sky130_fd_sc_hd__clkbuf_4 T4Y85__R0_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B574));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R0_INV_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9220));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R1_INV_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R2_INV_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R2_INV_1 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9256));
  sky130_fd_sc_hd__clkbuf_4 T4Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9292));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R0_INV_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y86__R1_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B583));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R1_INV_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R2_INV_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R2_INV_1 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9364));
  sky130_fd_sc_hd__clkbuf_4 T4Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9400));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R0_INV_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9436));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R1_INV_0 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R2_INV_0 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R2_INV_1 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y87__R3_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B37));
  sky130_fd_sc_hd__clkbuf_4 T4Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9508));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R0_INV_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9544));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R1_INV_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R2_INV_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R2_INV_1 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9580));
  sky130_fd_sc_hd__clkbuf_4 T4Y89__R0_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B601));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R0_INV_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9652));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R1_INV_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R2_INV_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R2_INV_1 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9688));
  sky130_fd_sc_hd__clkbuf_4 T4Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B869));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R0_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B905));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R1_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R2_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R2_INV_1 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B941));
  sky130_fd_sc_hd__clkbuf_4 T4Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B977));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R0_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1013));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R1_INV_0 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R2_INV_0 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R2_INV_1 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1049));
  sky130_fd_sc_hd__clkbuf_4 T5Y0__R0_BUF_0 (.A(clk_L1_B0), .X(clk_L0_B15));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R0_INV_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B50));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R1_INV_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R2_INV_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R2_INV_1 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B85));
  sky130_fd_sc_hd__clkbuf_4 T5Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1086));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R0_INV_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1122));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R1_INV_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R2_INV_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R2_INV_1 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1158));
  sky130_fd_sc_hd__clkbuf_4 T5Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1194));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R0_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1230));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R1_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R2_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R2_INV_1 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1266));
  sky130_fd_sc_hd__clkbuf_4 T5Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1302));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R0_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1338));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R1_INV_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R2_INV_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R2_INV_1 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1374));
  sky130_fd_sc_hd__clkbuf_4 T5Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1410));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R0_INV_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1446));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R1_INV_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R2_INV_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R2_INV_1 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1482));
  sky130_fd_sc_hd__clkbuf_4 T5Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1518));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R0_INV_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1553));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R1_INV_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R2_INV_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R2_INV_1 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1589));
  sky130_fd_sc_hd__clkbuf_4 T5Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1625));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R0_INV_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1661));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R1_INV_0 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R2_INV_0 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R2_INV_1 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1697));
  sky130_fd_sc_hd__clkbuf_4 T5Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1733));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R0_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1769));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R1_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R2_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R2_INV_1 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1805));
  sky130_fd_sc_hd__clkbuf_4 T5Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1841));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R0_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1877));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R1_INV_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R2_INV_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R2_INV_1 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1913));
  sky130_fd_sc_hd__clkbuf_4 T5Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1949));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R0_INV_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1985));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R1_INV_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R2_INV_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R2_INV_1 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2021));
  sky130_fd_sc_hd__clkbuf_4 T5Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2057));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R0_INV_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2093));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R1_INV_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R2_INV_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R2_INV_1 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2129));
  sky130_fd_sc_hd__clkbuf_4 T5Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B120));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R0_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B155));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R1_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R2_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R2_INV_1 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B190));
  sky130_fd_sc_hd__clkbuf_4 T5Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2165));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R0_INV_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2201));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R1_INV_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R2_INV_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R2_INV_1 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2237));
  sky130_fd_sc_hd__clkbuf_4 T5Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2273));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R0_INV_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2309));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R1_INV_0 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R2_INV_0 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R2_INV_1 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2345));
  sky130_fd_sc_hd__clkbuf_4 T5Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2381));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R0_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2417));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R1_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R2_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R2_INV_1 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2453));
  sky130_fd_sc_hd__clkbuf_4 T5Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2489));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R0_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2525));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R1_INV_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R2_INV_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R2_INV_1 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2561));
  sky130_fd_sc_hd__clkbuf_4 T5Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2597));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R0_INV_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2633));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R1_INV_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R2_INV_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R2_INV_1 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2669));
  sky130_fd_sc_hd__clkbuf_4 T5Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2705));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R0_INV_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2741));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R1_INV_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R2_INV_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R2_INV_1 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2777));
  sky130_fd_sc_hd__clkbuf_4 T5Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2813));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R0_INV_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2849));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R1_INV_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R2_INV_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R2_INV_1 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2885));
  sky130_fd_sc_hd__clkbuf_4 T5Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2921));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R0_INV_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2957));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R1_INV_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R2_INV_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R2_INV_1 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2993));
  sky130_fd_sc_hd__clkbuf_4 T5Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3029));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R0_INV_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3065));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R1_INV_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R2_INV_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R2_INV_1 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3101));
  sky130_fd_sc_hd__clkbuf_4 T5Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3137));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R0_INV_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3173));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R1_INV_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R2_INV_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R2_INV_1 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3209));
  sky130_fd_sc_hd__clkbuf_4 T5Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B225));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R0_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B260));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R1_INV_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R2_INV_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R2_INV_1 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B296));
  sky130_fd_sc_hd__clkbuf_4 T5Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3245));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R0_INV_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3281));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R1_INV_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R2_INV_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R2_INV_1 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3317));
  sky130_fd_sc_hd__clkbuf_4 T5Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3353));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R0_INV_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3389));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R1_INV_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R2_INV_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R2_INV_1 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3425));
  sky130_fd_sc_hd__clkbuf_4 T5Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3461));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R0_INV_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3497));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R1_INV_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R2_INV_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R2_INV_1 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3533));
  sky130_fd_sc_hd__clkbuf_4 T5Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3569));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R0_INV_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3605));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R1_INV_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R2_INV_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R2_INV_1 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3641));
  sky130_fd_sc_hd__clkbuf_4 T5Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3677));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R0_INV_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3713));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R1_INV_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R2_INV_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R2_INV_1 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3749));
  sky130_fd_sc_hd__clkbuf_4 T5Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3785));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R0_INV_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3821));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R1_INV_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R2_INV_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R2_INV_1 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3857));
  sky130_fd_sc_hd__clkbuf_4 T5Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3893));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R0_INV_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3929));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R1_INV_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R2_INV_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R2_INV_1 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3965));
  sky130_fd_sc_hd__clkbuf_4 T5Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4001));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R0_INV_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4037));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R1_INV_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R2_INV_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R2_INV_1 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4073));
  sky130_fd_sc_hd__clkbuf_4 T5Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4109));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R0_INV_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4145));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R1_INV_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R2_INV_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R2_INV_1 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4181));
  sky130_fd_sc_hd__clkbuf_4 T5Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4217));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R0_INV_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4253));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R1_INV_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R2_INV_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R2_INV_1 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4289));
  sky130_fd_sc_hd__clkbuf_4 T5Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B331));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R0_INV_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B366));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R1_INV_0 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R2_INV_0 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R2_INV_1 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B402));
  sky130_fd_sc_hd__clkbuf_4 T5Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4325));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R0_INV_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4361));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R1_INV_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R2_INV_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R2_INV_1 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4397));
  sky130_fd_sc_hd__clkbuf_4 T5Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4433));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R0_INV_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4469));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R1_INV_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R2_INV_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R2_INV_1 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4505));
  sky130_fd_sc_hd__clkbuf_4 T5Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4541));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R0_INV_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4577));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R1_INV_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R2_INV_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R2_INV_1 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4613));
  sky130_fd_sc_hd__clkbuf_4 T5Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4649));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R0_INV_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4685));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R1_INV_0 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R2_INV_0 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R2_INV_1 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4721));
  sky130_fd_sc_hd__clkbuf_4 T5Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4757));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R0_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4793));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R1_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R2_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R2_INV_1 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4829));
  sky130_fd_sc_hd__clkbuf_4 T5Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4865));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R0_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4901));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R1_INV_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R2_INV_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R2_INV_1 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4937));
  sky130_fd_sc_hd__clkbuf_4 T5Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4973));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R0_INV_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5009));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R1_INV_0 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R2_INV_0 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R2_INV_1 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5045));
  sky130_fd_sc_hd__clkbuf_4 T5Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5081));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R0_INV_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5117));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R1_INV_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R2_INV_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R2_INV_1 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5153));
  sky130_fd_sc_hd__clkbuf_4 T5Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5189));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R0_INV_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5225));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R1_INV_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R2_INV_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R2_INV_1 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5261));
  sky130_fd_sc_hd__clkbuf_4 T5Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5297));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R0_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5333));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R1_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R2_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R2_INV_1 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5369));
  sky130_fd_sc_hd__clkbuf_4 T5Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B438));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R0_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B474));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R1_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R2_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R2_INV_1 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B510));
  sky130_fd_sc_hd__clkbuf_4 T5Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5405));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R0_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5441));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R1_INV_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R2_INV_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R2_INV_1 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5477));
  sky130_fd_sc_hd__clkbuf_4 T5Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5513));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R0_INV_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5549));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R1_INV_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R2_INV_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R2_INV_1 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5585));
  sky130_fd_sc_hd__clkbuf_4 T5Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5621));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R0_INV_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5657));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R1_INV_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R2_INV_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R2_INV_1 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5693));
  sky130_fd_sc_hd__clkbuf_4 T5Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5729));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R0_INV_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5765));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R1_INV_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R2_INV_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R2_INV_1 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5801));
  sky130_fd_sc_hd__clkbuf_4 T5Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5837));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R0_INV_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5873));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R1_INV_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R2_INV_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R2_INV_1 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5909));
  sky130_fd_sc_hd__clkbuf_4 T5Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5945));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R0_INV_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5981));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R1_INV_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R2_INV_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R2_INV_1 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6017));
  sky130_fd_sc_hd__clkbuf_4 T5Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6053));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R0_INV_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6089));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R1_INV_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R2_INV_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R2_INV_1 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6125));
  sky130_fd_sc_hd__clkbuf_4 T5Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6161));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R0_INV_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6197));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R1_INV_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R2_INV_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R2_INV_1 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6233));
  sky130_fd_sc_hd__clkbuf_4 T5Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6269));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R0_INV_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6305));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R1_INV_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R2_INV_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R2_INV_1 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6341));
  sky130_fd_sc_hd__clkbuf_4 T5Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6377));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R0_INV_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6413));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R1_INV_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R2_INV_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R2_INV_1 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6449));
  sky130_fd_sc_hd__clkbuf_4 T5Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B546));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R0_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B582));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R1_INV_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R2_INV_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R2_INV_1 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B618));
  sky130_fd_sc_hd__clkbuf_4 T5Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6485));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R0_INV_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6521));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R1_INV_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R2_INV_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R2_INV_1 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6557));
  sky130_fd_sc_hd__clkbuf_4 T5Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6593));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R0_INV_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6629));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R1_INV_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R2_INV_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R2_INV_1 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6665));
  sky130_fd_sc_hd__clkbuf_4 T5Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6701));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R0_INV_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6737));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R1_INV_0 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R2_INV_0 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R2_INV_1 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6773));
  sky130_fd_sc_hd__clkbuf_4 T5Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6809));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R0_INV_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6845));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R1_INV_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R2_INV_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R2_INV_1 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6881));
  sky130_fd_sc_hd__clkbuf_4 T5Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6917));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R0_INV_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6953));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R1_INV_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R2_INV_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R2_INV_1 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6989));
  sky130_fd_sc_hd__clkbuf_4 T5Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7025));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R0_INV_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7061));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R1_INV_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R2_INV_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R2_INV_1 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7097));
  sky130_fd_sc_hd__clkbuf_4 T5Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7133));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R0_INV_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7169));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R1_INV_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R2_INV_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R2_INV_1 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7205));
  sky130_fd_sc_hd__clkbuf_4 T5Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7241));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R0_INV_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7277));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R1_INV_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R2_INV_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R2_INV_1 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7313));
  sky130_fd_sc_hd__clkbuf_4 T5Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7349));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R0_INV_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7385));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R1_INV_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R2_INV_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R2_INV_1 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7421));
  sky130_fd_sc_hd__clkbuf_4 T5Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7457));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R0_INV_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7493));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R1_INV_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R2_INV_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R2_INV_1 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7529));
  sky130_fd_sc_hd__clkbuf_4 T5Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B654));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R0_INV_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B690));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R1_INV_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R2_INV_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R2_INV_1 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B726));
  sky130_fd_sc_hd__clkbuf_4 T5Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7565));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R0_INV_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7601));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R1_INV_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R2_INV_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R2_INV_1 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7637));
  sky130_fd_sc_hd__clkbuf_4 T5Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7673));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R0_INV_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7709));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R1_INV_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R2_INV_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R2_INV_1 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7745));
  sky130_fd_sc_hd__clkbuf_4 T5Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7781));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R0_INV_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7817));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R1_INV_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R2_INV_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R2_INV_1 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7853));
  sky130_fd_sc_hd__clkbuf_4 T5Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7889));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R0_INV_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7925));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R1_INV_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R2_INV_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R2_INV_1 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7961));
  sky130_fd_sc_hd__clkbuf_4 T5Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7997));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R0_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8033));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R1_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R2_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R2_INV_1 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8069));
  sky130_fd_sc_hd__clkbuf_4 T5Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8105));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R0_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8141));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R1_INV_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R2_INV_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R2_INV_1 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8177));
  sky130_fd_sc_hd__clkbuf_4 T5Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8213));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R0_INV_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8249));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R1_INV_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R2_INV_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R2_INV_1 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8285));
  sky130_fd_sc_hd__clkbuf_4 T5Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8321));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R0_INV_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8357));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R1_INV_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R2_INV_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R2_INV_1 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8393));
  sky130_fd_sc_hd__clkbuf_4 T5Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8429));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R0_INV_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8465));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R1_INV_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R2_INV_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R2_INV_1 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8501));
  sky130_fd_sc_hd__clkbuf_4 T5Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8537));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R0_INV_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8573));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R1_INV_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R2_INV_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R2_INV_1 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8609));
  sky130_fd_sc_hd__clkbuf_4 T5Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B762));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R0_INV_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B798));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R1_INV_0 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R2_INV_0 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R2_INV_1 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B834));
  sky130_fd_sc_hd__clkbuf_4 T5Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8645));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R0_INV_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8681));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R1_INV_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R2_INV_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R2_INV_1 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8717));
  sky130_fd_sc_hd__clkbuf_4 T5Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8753));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R0_INV_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8789));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R1_INV_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R2_INV_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R2_INV_1 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8825));
  sky130_fd_sc_hd__clkbuf_4 T5Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8861));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R0_INV_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8897));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R1_INV_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R2_INV_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R2_INV_1 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8933));
  sky130_fd_sc_hd__clkbuf_4 T5Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8969));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R0_INV_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9005));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R1_INV_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R2_INV_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R2_INV_1 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9041));
  sky130_fd_sc_hd__clkbuf_4 T5Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9077));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R0_INV_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9113));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R1_INV_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R2_INV_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R2_INV_1 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9149));
  sky130_fd_sc_hd__clkbuf_4 T5Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9185));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R0_INV_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9221));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R1_INV_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R2_INV_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R2_INV_1 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9257));
  sky130_fd_sc_hd__clkbuf_4 T5Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9293));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R0_INV_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9329));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R1_INV_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R2_INV_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R2_INV_1 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9365));
  sky130_fd_sc_hd__clkbuf_4 T5Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9401));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R0_INV_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9437));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R1_INV_0 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R2_INV_0 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R2_INV_1 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9473));
  sky130_fd_sc_hd__clkbuf_4 T5Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9509));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R0_INV_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9545));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R1_INV_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R2_INV_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R2_INV_1 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9581));
  sky130_fd_sc_hd__clkbuf_4 T5Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9617));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R0_INV_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9653));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R1_INV_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R2_INV_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R2_INV_1 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9689));
  sky130_fd_sc_hd__clkbuf_4 T5Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B870));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R0_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B906));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R1_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R2_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R2_INV_1 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B942));
  sky130_fd_sc_hd__clkbuf_4 T5Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B978));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R0_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1014));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R1_INV_0 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R2_INV_0 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R2_INV_1 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1050));
  sky130_fd_sc_hd__clkbuf_4 T6Y0__R0_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B1));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R0_INV_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B51));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R1_INV_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R2_INV_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R2_INV_1 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B86));
  sky130_fd_sc_hd__clkbuf_4 T6Y10__R0_BUF_0 (.A(clk_L1_B67), .X(clk_L0_B1087));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R0_INV_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1123));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R1_INV_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R2_INV_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R2_INV_1 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1159));
  sky130_fd_sc_hd__clkbuf_4 T6Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1195));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R0_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y11__R1_BUF_0 (.A(clk_L1_B76), .X(clk_L0_B1231));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R1_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R2_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R2_INV_1 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1267));
  sky130_fd_sc_hd__clkbuf_4 T6Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1303));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R0_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1339));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R1_INV_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R2_INV_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R2_INV_1 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y12__R3_BUF_0 (.A(clk_L1_B85), .X(clk_L0_B1375));
  sky130_fd_sc_hd__clkbuf_4 T6Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1411));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R0_INV_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1447));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R1_INV_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R2_INV_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R2_INV_1 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1483));
  sky130_fd_sc_hd__clkbuf_4 T6Y14__R0_BUF_0 (.A(clk_L1_B94), .X(clk_L0_B1519));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R0_INV_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1554));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R1_INV_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R2_INV_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R2_INV_1 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1590));
  sky130_fd_sc_hd__clkbuf_4 T6Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1626));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R0_INV_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1662));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R1_INV_0 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R2_INV_0 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R2_INV_1 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1698));
  sky130_fd_sc_hd__clkbuf_4 T6Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1734));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R0_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1770));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R1_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R2_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R2_INV_1 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1806));
  sky130_fd_sc_hd__clkbuf_4 T6Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1842));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R0_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1878));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R1_INV_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R2_INV_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R2_INV_1 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1914));
  sky130_fd_sc_hd__clkbuf_4 T6Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1950));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R0_INV_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1986));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R1_INV_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R2_INV_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R2_INV_1 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2022));
  sky130_fd_sc_hd__clkbuf_4 T6Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2058));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R0_INV_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2094));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R1_INV_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R2_INV_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R2_INV_1 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2130));
  sky130_fd_sc_hd__clkbuf_4 T6Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B121));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R0_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B156));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R1_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R2_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R2_INV_1 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y1__R3_BUF_0 (.A(clk_L1_B11), .X(clk_L0_B191));
  sky130_fd_sc_hd__clkbuf_4 T6Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2166));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R0_INV_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2202));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R1_INV_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R2_INV_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R2_INV_1 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2238));
  sky130_fd_sc_hd__clkbuf_4 T6Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2274));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R0_INV_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2310));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R1_INV_0 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R2_INV_0 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R2_INV_1 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2346));
  sky130_fd_sc_hd__clkbuf_4 T6Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2382));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R0_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2418));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R1_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R2_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R2_INV_1 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2454));
  sky130_fd_sc_hd__clkbuf_4 T6Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2490));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R0_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2526));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R1_INV_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R2_INV_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R2_INV_1 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2562));
  sky130_fd_sc_hd__clkbuf_4 T6Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2598));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R0_INV_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2634));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R1_INV_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R2_INV_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R2_INV_1 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2670));
  sky130_fd_sc_hd__clkbuf_4 T6Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2706));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R0_INV_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2742));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R1_INV_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R2_INV_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R2_INV_1 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2778));
  sky130_fd_sc_hd__clkbuf_4 T6Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2814));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R0_INV_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2850));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R1_INV_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R2_INV_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R2_INV_1 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2886));
  sky130_fd_sc_hd__clkbuf_4 T6Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2922));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R0_INV_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2958));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R1_INV_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R2_INV_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R2_INV_1 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2994));
  sky130_fd_sc_hd__clkbuf_4 T6Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3030));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R0_INV_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3066));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R1_INV_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R2_INV_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R2_INV_1 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3102));
  sky130_fd_sc_hd__clkbuf_4 T6Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3138));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R0_INV_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3174));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R1_INV_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R2_INV_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R2_INV_1 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3210));
  sky130_fd_sc_hd__clkbuf_4 T6Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B226));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R0_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B261));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R1_INV_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R2_INV_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R2_INV_1 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B297));
  sky130_fd_sc_hd__clkbuf_4 T6Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3246));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R0_INV_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3282));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R1_INV_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R2_INV_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R2_INV_1 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3318));
  sky130_fd_sc_hd__clkbuf_4 T6Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3354));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R0_INV_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3390));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R1_INV_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R2_INV_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R2_INV_1 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3426));
  sky130_fd_sc_hd__clkbuf_4 T6Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3462));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R0_INV_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3498));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R1_INV_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R2_INV_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R2_INV_1 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3534));
  sky130_fd_sc_hd__clkbuf_4 T6Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3570));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R0_INV_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3606));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R1_INV_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R2_INV_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R2_INV_1 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3642));
  sky130_fd_sc_hd__clkbuf_4 T6Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3678));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R0_INV_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3714));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R1_INV_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R2_INV_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R2_INV_1 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3750));
  sky130_fd_sc_hd__clkbuf_4 T6Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3786));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R0_INV_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3822));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R1_INV_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R2_INV_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R2_INV_1 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3858));
  sky130_fd_sc_hd__clkbuf_4 T6Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3894));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R0_INV_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3930));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R1_INV_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R2_INV_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R2_INV_1 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3966));
  sky130_fd_sc_hd__clkbuf_4 T6Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4002));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R0_INV_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4038));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R1_INV_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R2_INV_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R2_INV_1 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4074));
  sky130_fd_sc_hd__clkbuf_4 T6Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4110));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R0_INV_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4146));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R1_INV_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R2_INV_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R2_INV_1 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4182));
  sky130_fd_sc_hd__clkbuf_4 T6Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4218));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R0_INV_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4254));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R1_INV_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R2_INV_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R2_INV_1 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4290));
  sky130_fd_sc_hd__clkbuf_4 T6Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B332));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R0_INV_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y3__R1_BUF_0 (.A(clk_L1_B22), .X(clk_L0_B367));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R1_INV_0 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R2_INV_0 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R2_INV_1 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B403));
  sky130_fd_sc_hd__clkbuf_4 T6Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4326));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R0_INV_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4362));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R1_INV_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R2_INV_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R2_INV_1 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4398));
  sky130_fd_sc_hd__clkbuf_4 T6Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4434));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R0_INV_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4470));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R1_INV_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R2_INV_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R2_INV_1 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4506));
  sky130_fd_sc_hd__clkbuf_4 T6Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4542));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R0_INV_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4578));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R1_INV_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R2_INV_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R2_INV_1 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4614));
  sky130_fd_sc_hd__clkbuf_4 T6Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4650));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R0_INV_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4686));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R1_INV_0 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R2_INV_0 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R2_INV_1 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4722));
  sky130_fd_sc_hd__clkbuf_4 T6Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4758));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R0_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4794));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R1_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R2_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R2_INV_1 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4830));
  sky130_fd_sc_hd__clkbuf_4 T6Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4866));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R0_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4902));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R1_INV_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R2_INV_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R2_INV_1 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4938));
  sky130_fd_sc_hd__clkbuf_4 T6Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4974));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R0_INV_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5010));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R1_INV_0 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R2_INV_0 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R2_INV_1 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5046));
  sky130_fd_sc_hd__clkbuf_4 T6Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5082));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R0_INV_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5118));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R1_INV_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R2_INV_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R2_INV_1 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5154));
  sky130_fd_sc_hd__clkbuf_4 T6Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5190));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R0_INV_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5226));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R1_INV_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R2_INV_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R2_INV_1 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5262));
  sky130_fd_sc_hd__clkbuf_4 T6Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5298));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R0_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5334));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R1_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R2_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R2_INV_1 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5370));
  sky130_fd_sc_hd__clkbuf_4 T6Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B439));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R0_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B475));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R1_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R2_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R2_INV_1 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y4__R3_BUF_0 (.A(clk_L1_B31), .X(clk_L0_B511));
  sky130_fd_sc_hd__clkbuf_4 T6Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5406));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R0_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5442));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R1_INV_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R2_INV_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R2_INV_1 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5478));
  sky130_fd_sc_hd__clkbuf_4 T6Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5514));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R0_INV_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5550));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R1_INV_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R2_INV_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R2_INV_1 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5586));
  sky130_fd_sc_hd__clkbuf_4 T6Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5622));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R0_INV_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5658));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R1_INV_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R2_INV_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R2_INV_1 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5694));
  sky130_fd_sc_hd__clkbuf_4 T6Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5730));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R0_INV_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5766));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R1_INV_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R2_INV_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R2_INV_1 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5802));
  sky130_fd_sc_hd__clkbuf_4 T6Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5838));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R0_INV_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5874));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R1_INV_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R2_INV_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R2_INV_1 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5910));
  sky130_fd_sc_hd__clkbuf_4 T6Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5946));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R0_INV_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5982));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R1_INV_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R2_INV_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R2_INV_1 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6018));
  sky130_fd_sc_hd__clkbuf_4 T6Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6054));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R0_INV_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6090));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R1_INV_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R2_INV_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R2_INV_1 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6126));
  sky130_fd_sc_hd__clkbuf_4 T6Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6162));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R0_INV_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6198));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R1_INV_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R2_INV_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R2_INV_1 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6234));
  sky130_fd_sc_hd__clkbuf_4 T6Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6270));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R0_INV_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6306));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R1_INV_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R2_INV_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R2_INV_1 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6342));
  sky130_fd_sc_hd__clkbuf_4 T6Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6378));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R0_INV_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6414));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R1_INV_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R2_INV_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R2_INV_1 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6450));
  sky130_fd_sc_hd__clkbuf_4 T6Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B547));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R0_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B583));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R1_INV_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R2_INV_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R2_INV_1 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B619));
  sky130_fd_sc_hd__clkbuf_4 T6Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6486));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R0_INV_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6522));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R1_INV_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R2_INV_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R2_INV_1 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6558));
  sky130_fd_sc_hd__clkbuf_4 T6Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6594));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R0_INV_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6630));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R1_INV_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R2_INV_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R2_INV_1 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6666));
  sky130_fd_sc_hd__clkbuf_4 T6Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6702));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R0_INV_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6738));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R1_INV_0 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R2_INV_0 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R2_INV_1 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6774));
  sky130_fd_sc_hd__clkbuf_4 T6Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6810));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R0_INV_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6846));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R1_INV_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R2_INV_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R2_INV_1 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6882));
  sky130_fd_sc_hd__clkbuf_4 T6Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6918));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R0_INV_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6954));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R1_INV_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R2_INV_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R2_INV_1 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6990));
  sky130_fd_sc_hd__clkbuf_4 T6Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7026));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R0_INV_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7062));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R1_INV_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R2_INV_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R2_INV_1 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7098));
  sky130_fd_sc_hd__clkbuf_4 T6Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7134));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R0_INV_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7170));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R1_INV_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R2_INV_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R2_INV_1 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7206));
  sky130_fd_sc_hd__clkbuf_4 T6Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7242));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R0_INV_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7278));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R1_INV_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R2_INV_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R2_INV_1 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7314));
  sky130_fd_sc_hd__clkbuf_4 T6Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7350));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R0_INV_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7386));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R1_INV_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R2_INV_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R2_INV_1 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7422));
  sky130_fd_sc_hd__clkbuf_4 T6Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7458));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R0_INV_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7494));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R1_INV_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R2_INV_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R2_INV_1 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7530));
  sky130_fd_sc_hd__clkbuf_4 T6Y6__R0_BUF_0 (.A(clk_L1_B40), .X(clk_L0_B655));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R0_INV_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B691));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R1_INV_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R2_INV_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R2_INV_1 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B727));
  sky130_fd_sc_hd__clkbuf_4 T6Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7566));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R0_INV_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7602));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R1_INV_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R2_INV_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R2_INV_1 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7638));
  sky130_fd_sc_hd__clkbuf_4 T6Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7674));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R0_INV_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7710));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R1_INV_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R2_INV_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R2_INV_1 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7746));
  sky130_fd_sc_hd__clkbuf_4 T6Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7782));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R0_INV_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7818));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R1_INV_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R2_INV_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R2_INV_1 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7854));
  sky130_fd_sc_hd__clkbuf_4 T6Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7890));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R0_INV_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7926));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R1_INV_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R2_INV_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R2_INV_1 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7962));
  sky130_fd_sc_hd__clkbuf_4 T6Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7998));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R0_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8034));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R1_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R2_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R2_INV_1 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8070));
  sky130_fd_sc_hd__clkbuf_4 T6Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8106));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R0_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8142));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R1_INV_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R2_INV_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R2_INV_1 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8178));
  sky130_fd_sc_hd__clkbuf_4 T6Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8214));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R0_INV_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8250));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R1_INV_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R2_INV_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R2_INV_1 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8286));
  sky130_fd_sc_hd__clkbuf_4 T6Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8322));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R0_INV_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8358));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R1_INV_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R2_INV_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R2_INV_1 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8394));
  sky130_fd_sc_hd__clkbuf_4 T6Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8430));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R0_INV_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8466));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R1_INV_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R2_INV_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R2_INV_1 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8502));
  sky130_fd_sc_hd__clkbuf_4 T6Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8538));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R0_INV_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8574));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R1_INV_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R2_INV_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R2_INV_1 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8610));
  sky130_fd_sc_hd__clkbuf_4 T6Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B763));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R0_INV_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y7__R1_BUF_0 (.A(clk_L1_B49), .X(clk_L0_B799));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R1_INV_0 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R2_INV_0 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R2_INV_1 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B835));
  sky130_fd_sc_hd__clkbuf_4 T6Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8646));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R0_INV_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8682));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R1_INV_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R2_INV_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R2_INV_1 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8718));
  sky130_fd_sc_hd__clkbuf_4 T6Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8754));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R0_INV_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8790));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R1_INV_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R2_INV_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R2_INV_1 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8826));
  sky130_fd_sc_hd__clkbuf_4 T6Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8862));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R0_INV_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8898));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R1_INV_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R2_INV_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R2_INV_1 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8934));
  sky130_fd_sc_hd__clkbuf_4 T6Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8970));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R0_INV_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9006));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R1_INV_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R2_INV_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R2_INV_1 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9042));
  sky130_fd_sc_hd__clkbuf_4 T6Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9078));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R0_INV_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9114));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R1_INV_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R2_INV_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R2_INV_1 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9150));
  sky130_fd_sc_hd__clkbuf_4 T6Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9186));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R0_INV_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9222));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R1_INV_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R2_INV_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R2_INV_1 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9258));
  sky130_fd_sc_hd__clkbuf_4 T6Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9294));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R0_INV_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9330));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R1_INV_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R2_INV_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R2_INV_1 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9366));
  sky130_fd_sc_hd__clkbuf_4 T6Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9402));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R0_INV_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9438));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R1_INV_0 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R2_INV_0 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R2_INV_1 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9474));
  sky130_fd_sc_hd__clkbuf_4 T6Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9510));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R0_INV_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9546));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R1_INV_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R2_INV_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R2_INV_1 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9582));
  sky130_fd_sc_hd__clkbuf_4 T6Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9618));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R0_INV_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9654));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R1_INV_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R2_INV_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R2_INV_1 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9690));
  sky130_fd_sc_hd__clkbuf_4 T6Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B871));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R0_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B907));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R1_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R2_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R2_INV_1 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y8__R3_BUF_0 (.A(clk_L1_B58), .X(clk_L0_B943));
  sky130_fd_sc_hd__clkbuf_4 T6Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B979));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R0_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1015));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R1_INV_0 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R2_INV_0 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R2_INV_1 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1051));
  sky130_fd_sc_hd__clkbuf_4 T7Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B17));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R0_INV_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B52));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R1_INV_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R2_INV_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R2_INV_1 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B87));
  sky130_fd_sc_hd__clkbuf_4 T7Y10__R0_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B68));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R0_INV_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1124));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R1_INV_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R2_INV_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R2_INV_1 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1160));
  sky130_fd_sc_hd__clkbuf_4 T7Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1196));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R0_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y11__R1_BUF_0 (.A(clk_L2_B4), .X(clk_L1_B77));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R1_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R2_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R2_INV_1 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1268));
  sky130_fd_sc_hd__clkbuf_4 T7Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1304));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R0_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1340));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R1_INV_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R2_INV_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R2_INV_1 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y12__R3_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B86));
  sky130_fd_sc_hd__clkbuf_4 T7Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1412));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R0_INV_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1448));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R1_INV_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R2_INV_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R2_INV_1 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1484));
  sky130_fd_sc_hd__clkbuf_4 T7Y14__R0_BUF_0 (.A(clk_L2_B5), .X(clk_L1_B95));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R0_INV_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1555));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R1_INV_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R2_INV_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R2_INV_1 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1591));
  sky130_fd_sc_hd__clkbuf_4 T7Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1627));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R0_INV_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y15__R1_BUF_0 (.A(clk_L1_B103), .X(clk_L0_B1663));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R1_INV_0 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R2_INV_0 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R2_INV_1 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1699));
  sky130_fd_sc_hd__clkbuf_4 T7Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1735));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R0_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1771));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R1_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R2_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R2_INV_1 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y16__R3_BUF_0 (.A(clk_L1_B112), .X(clk_L0_B1807));
  sky130_fd_sc_hd__clkbuf_4 T7Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1843));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R0_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1879));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R1_INV_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R2_INV_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R2_INV_1 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1915));
  sky130_fd_sc_hd__clkbuf_4 T7Y18__R0_BUF_0 (.A(clk_L1_B121), .X(clk_L0_B1951));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R0_INV_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1987));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R1_INV_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R2_INV_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R2_INV_1 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2023));
  sky130_fd_sc_hd__clkbuf_4 T7Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2059));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R0_INV_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y19__R1_BUF_0 (.A(clk_L1_B130), .X(clk_L0_B2095));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R1_INV_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R2_INV_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R2_INV_1 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2131));
  sky130_fd_sc_hd__clkbuf_4 T7Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B122));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R0_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B157));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R1_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R2_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R2_INV_1 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y1__R3_BUF_0 (.A(clk_L2_B0), .X(clk_L1_B12));
  sky130_fd_sc_hd__clkbuf_4 T7Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2167));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R0_INV_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2203));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R1_INV_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R2_INV_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R2_INV_1 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y20__R3_BUF_0 (.A(clk_L1_B139), .X(clk_L0_B2239));
  sky130_fd_sc_hd__clkbuf_4 T7Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2275));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R0_INV_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2311));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R1_INV_0 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R2_INV_0 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R2_INV_1 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2347));
  sky130_fd_sc_hd__clkbuf_4 T7Y22__R0_BUF_0 (.A(clk_L1_B148), .X(clk_L0_B2383));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R0_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2419));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R1_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R2_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R2_INV_1 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2455));
  sky130_fd_sc_hd__clkbuf_4 T7Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2491));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R0_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y23__R1_BUF_0 (.A(clk_L1_B157), .X(clk_L0_B2527));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R1_INV_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R2_INV_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R2_INV_1 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2563));
  sky130_fd_sc_hd__clkbuf_4 T7Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2599));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R0_INV_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2635));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R1_INV_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R2_INV_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R2_INV_1 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y24__R3_BUF_0 (.A(clk_L1_B166), .X(clk_L0_B2671));
  sky130_fd_sc_hd__clkbuf_4 T7Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2707));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R0_INV_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2743));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R1_INV_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R2_INV_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R2_INV_1 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2779));
  sky130_fd_sc_hd__clkbuf_4 T7Y26__R0_BUF_0 (.A(clk_L1_B175), .X(clk_L0_B2815));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R0_INV_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2851));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R1_INV_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R2_INV_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R2_INV_1 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2887));
  sky130_fd_sc_hd__clkbuf_4 T7Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2923));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R0_INV_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y27__R1_BUF_0 (.A(clk_L1_B184), .X(clk_L0_B2959));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R1_INV_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R2_INV_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R2_INV_1 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2995));
  sky130_fd_sc_hd__clkbuf_4 T7Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3031));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R0_INV_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3067));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R1_INV_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R2_INV_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R2_INV_1 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y28__R3_BUF_0 (.A(clk_L1_B193), .X(clk_L0_B3103));
  sky130_fd_sc_hd__clkbuf_4 T7Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3139));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R0_INV_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3175));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R1_INV_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R2_INV_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R2_INV_1 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3211));
  sky130_fd_sc_hd__clkbuf_4 T7Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B227));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R0_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B262));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R1_INV_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R2_INV_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R2_INV_1 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B298));
  sky130_fd_sc_hd__clkbuf_4 T7Y30__R0_BUF_0 (.A(clk_L1_B202), .X(clk_L0_B3247));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R0_INV_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3283));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R1_INV_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R2_INV_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R2_INV_1 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3319));
  sky130_fd_sc_hd__clkbuf_4 T7Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3355));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R0_INV_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y31__R1_BUF_0 (.A(clk_L1_B211), .X(clk_L0_B3391));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R1_INV_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R2_INV_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R2_INV_1 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3427));
  sky130_fd_sc_hd__clkbuf_4 T7Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3463));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R0_INV_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3499));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R1_INV_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R2_INV_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R2_INV_1 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y32__R3_BUF_0 (.A(clk_L1_B220), .X(clk_L0_B3535));
  sky130_fd_sc_hd__clkbuf_4 T7Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3571));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R0_INV_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3607));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R1_INV_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R2_INV_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R2_INV_1 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3643));
  sky130_fd_sc_hd__clkbuf_4 T7Y34__R0_BUF_0 (.A(clk_L1_B229), .X(clk_L0_B3679));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R0_INV_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3715));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R1_INV_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R2_INV_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R2_INV_1 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3751));
  sky130_fd_sc_hd__clkbuf_4 T7Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3787));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R0_INV_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y35__R1_BUF_0 (.A(clk_L1_B238), .X(clk_L0_B3823));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R1_INV_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R2_INV_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R2_INV_1 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3859));
  sky130_fd_sc_hd__clkbuf_4 T7Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3895));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R0_INV_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3931));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R1_INV_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R2_INV_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R2_INV_1 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y36__R3_BUF_0 (.A(clk_L1_B247), .X(clk_L0_B3967));
  sky130_fd_sc_hd__clkbuf_4 T7Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4003));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R0_INV_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4039));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R1_INV_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R2_INV_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R2_INV_1 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4075));
  sky130_fd_sc_hd__clkbuf_4 T7Y38__R0_BUF_0 (.A(clk_L1_B256), .X(clk_L0_B4111));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R0_INV_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4147));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R1_INV_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R2_INV_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R2_INV_1 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4183));
  sky130_fd_sc_hd__clkbuf_4 T7Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4219));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R0_INV_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y39__R1_BUF_0 (.A(clk_L1_B265), .X(clk_L0_B4255));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R1_INV_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R2_INV_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R2_INV_1 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4291));
  sky130_fd_sc_hd__clkbuf_4 T7Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B333));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R0_INV_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y3__R1_BUF_0 (.A(clk_L2_B1), .X(clk_L1_B23));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R1_INV_0 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R2_INV_0 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R2_INV_1 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B404));
  sky130_fd_sc_hd__clkbuf_4 T7Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4327));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R0_INV_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4363));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R1_INV_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R2_INV_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R2_INV_1 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y40__R3_BUF_0 (.A(clk_L1_B274), .X(clk_L0_B4399));
  sky130_fd_sc_hd__clkbuf_4 T7Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4435));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R0_INV_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4471));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R1_INV_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R2_INV_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R2_INV_1 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4507));
  sky130_fd_sc_hd__clkbuf_4 T7Y42__R0_BUF_0 (.A(clk_L1_B283), .X(clk_L0_B4543));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R0_INV_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4579));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R1_INV_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R2_INV_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R2_INV_1 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4615));
  sky130_fd_sc_hd__clkbuf_4 T7Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4651));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R0_INV_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y43__R1_BUF_0 (.A(clk_L1_B292), .X(clk_L0_B4687));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R1_INV_0 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R2_INV_0 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R2_INV_1 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4723));
  sky130_fd_sc_hd__clkbuf_4 T7Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4759));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R0_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4795));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R1_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R2_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R2_INV_1 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y44__R3_BUF_0 (.A(clk_L1_B301), .X(clk_L0_B4831));
  sky130_fd_sc_hd__clkbuf_4 T7Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4867));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R0_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4903));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R1_INV_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R2_INV_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R2_INV_1 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4939));
  sky130_fd_sc_hd__clkbuf_4 T7Y46__R0_BUF_0 (.A(clk_L1_B310), .X(clk_L0_B4975));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R0_INV_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5011));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R1_INV_0 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R2_INV_0 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R2_INV_1 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5047));
  sky130_fd_sc_hd__clkbuf_4 T7Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5083));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R0_INV_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y47__R1_BUF_0 (.A(clk_L1_B319), .X(clk_L0_B5119));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R1_INV_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R2_INV_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R2_INV_1 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5155));
  sky130_fd_sc_hd__clkbuf_4 T7Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5191));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R0_INV_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5227));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R1_INV_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R2_INV_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R2_INV_1 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y48__R3_BUF_0 (.A(clk_L1_B328), .X(clk_L0_B5263));
  sky130_fd_sc_hd__clkbuf_4 T7Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5299));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R0_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5335));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R1_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R2_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R2_INV_1 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5371));
  sky130_fd_sc_hd__clkbuf_4 T7Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B440));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R0_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B476));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R1_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R2_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R2_INV_1 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y4__R3_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B2));
  sky130_fd_sc_hd__clkbuf_4 T7Y50__R0_BUF_0 (.A(clk_L1_B337), .X(clk_L0_B5407));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R0_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5443));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R1_INV_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R2_INV_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R2_INV_1 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5479));
  sky130_fd_sc_hd__clkbuf_4 T7Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5515));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R0_INV_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y51__R1_BUF_0 (.A(clk_L1_B346), .X(clk_L0_B5551));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R1_INV_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R2_INV_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R2_INV_1 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5587));
  sky130_fd_sc_hd__clkbuf_4 T7Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5623));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R0_INV_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5659));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R1_INV_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R2_INV_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R2_INV_1 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y52__R3_BUF_0 (.A(clk_L1_B355), .X(clk_L0_B5695));
  sky130_fd_sc_hd__clkbuf_4 T7Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5731));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R0_INV_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5767));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R1_INV_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R2_INV_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R2_INV_1 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5803));
  sky130_fd_sc_hd__clkbuf_4 T7Y54__R0_BUF_0 (.A(clk_L1_B364), .X(clk_L0_B5839));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R0_INV_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5875));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R1_INV_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R2_INV_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R2_INV_1 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5911));
  sky130_fd_sc_hd__clkbuf_4 T7Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5947));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R0_INV_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y55__R1_BUF_0 (.A(clk_L1_B373), .X(clk_L0_B5983));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R1_INV_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R2_INV_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R2_INV_1 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6019));
  sky130_fd_sc_hd__clkbuf_4 T7Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6055));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R0_INV_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6091));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R1_INV_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R2_INV_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R2_INV_1 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y56__R3_BUF_0 (.A(clk_L1_B382), .X(clk_L0_B6127));
  sky130_fd_sc_hd__clkbuf_4 T7Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6163));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R0_INV_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6199));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R1_INV_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R2_INV_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R2_INV_1 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6235));
  sky130_fd_sc_hd__clkbuf_4 T7Y58__R0_BUF_0 (.A(clk_L1_B391), .X(clk_L0_B6271));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R0_INV_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6307));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R1_INV_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R2_INV_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R2_INV_1 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6343));
  sky130_fd_sc_hd__clkbuf_4 T7Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6379));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R0_INV_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y59__R1_BUF_0 (.A(clk_L1_B400), .X(clk_L0_B6415));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R1_INV_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R2_INV_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R2_INV_1 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6451));
  sky130_fd_sc_hd__clkbuf_4 T7Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B548));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R0_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B584));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R1_INV_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R2_INV_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R2_INV_1 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B620));
  sky130_fd_sc_hd__clkbuf_4 T7Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6487));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R0_INV_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6523));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R1_INV_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R2_INV_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R2_INV_1 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y60__R3_BUF_0 (.A(clk_L1_B409), .X(clk_L0_B6559));
  sky130_fd_sc_hd__clkbuf_4 T7Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6595));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R0_INV_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6631));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R1_INV_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R2_INV_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R2_INV_1 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6667));
  sky130_fd_sc_hd__clkbuf_4 T7Y62__R0_BUF_0 (.A(clk_L1_B418), .X(clk_L0_B6703));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R0_INV_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6739));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R1_INV_0 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R2_INV_0 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R2_INV_1 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6775));
  sky130_fd_sc_hd__clkbuf_4 T7Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6811));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R0_INV_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y63__R1_BUF_0 (.A(clk_L1_B427), .X(clk_L0_B6847));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R1_INV_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R2_INV_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R2_INV_1 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6883));
  sky130_fd_sc_hd__clkbuf_4 T7Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6919));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R0_INV_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6955));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R1_INV_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R2_INV_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R2_INV_1 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y64__R3_BUF_0 (.A(clk_L1_B436), .X(clk_L0_B6991));
  sky130_fd_sc_hd__clkbuf_4 T7Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7027));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R0_INV_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7063));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R1_INV_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R2_INV_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R2_INV_1 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7099));
  sky130_fd_sc_hd__clkbuf_4 T7Y66__R0_BUF_0 (.A(clk_L1_B445), .X(clk_L0_B7135));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R0_INV_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7171));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R1_INV_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R2_INV_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R2_INV_1 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7207));
  sky130_fd_sc_hd__clkbuf_4 T7Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7243));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R0_INV_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y67__R1_BUF_0 (.A(clk_L1_B454), .X(clk_L0_B7279));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R1_INV_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R2_INV_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R2_INV_1 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7315));
  sky130_fd_sc_hd__clkbuf_4 T7Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7351));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R0_INV_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7387));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R1_INV_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R2_INV_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R2_INV_1 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y68__R3_BUF_0 (.A(clk_L1_B463), .X(clk_L0_B7423));
  sky130_fd_sc_hd__clkbuf_4 T7Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7459));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R0_INV_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7495));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R1_INV_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R2_INV_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R2_INV_1 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7531));
  sky130_fd_sc_hd__clkbuf_4 T7Y6__R0_BUF_0 (.A(clk_L2_B2), .X(clk_L1_B41));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R0_INV_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B692));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R1_INV_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R2_INV_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R2_INV_1 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B728));
  sky130_fd_sc_hd__clkbuf_4 T7Y70__R0_BUF_0 (.A(clk_L1_B472), .X(clk_L0_B7567));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R0_INV_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7603));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R1_INV_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R2_INV_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R2_INV_1 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7639));
  sky130_fd_sc_hd__clkbuf_4 T7Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7675));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R0_INV_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y71__R1_BUF_0 (.A(clk_L1_B481), .X(clk_L0_B7711));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R1_INV_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R2_INV_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R2_INV_1 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7747));
  sky130_fd_sc_hd__clkbuf_4 T7Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7783));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R0_INV_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7819));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R1_INV_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R2_INV_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R2_INV_1 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y72__R3_BUF_0 (.A(clk_L1_B490), .X(clk_L0_B7855));
  sky130_fd_sc_hd__clkbuf_4 T7Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7891));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R0_INV_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7927));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R1_INV_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R2_INV_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R2_INV_1 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7963));
  sky130_fd_sc_hd__clkbuf_4 T7Y74__R0_BUF_0 (.A(clk_L1_B499), .X(clk_L0_B7999));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R0_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8035));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R1_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R2_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R2_INV_1 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8071));
  sky130_fd_sc_hd__clkbuf_4 T7Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8107));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R0_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y75__R1_BUF_0 (.A(clk_L1_B508), .X(clk_L0_B8143));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R1_INV_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R2_INV_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R2_INV_1 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8179));
  sky130_fd_sc_hd__clkbuf_4 T7Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8215));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R0_INV_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8251));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R1_INV_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R2_INV_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R2_INV_1 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y76__R3_BUF_0 (.A(clk_L1_B517), .X(clk_L0_B8287));
  sky130_fd_sc_hd__clkbuf_4 T7Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8323));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R0_INV_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8359));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R1_INV_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R2_INV_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R2_INV_1 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8395));
  sky130_fd_sc_hd__clkbuf_4 T7Y78__R0_BUF_0 (.A(clk_L1_B526), .X(clk_L0_B8431));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R0_INV_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8467));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R1_INV_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R2_INV_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R2_INV_1 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8503));
  sky130_fd_sc_hd__clkbuf_4 T7Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8539));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R0_INV_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y79__R1_BUF_0 (.A(clk_L1_B535), .X(clk_L0_B8575));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R1_INV_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R2_INV_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R2_INV_1 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8611));
  sky130_fd_sc_hd__clkbuf_4 T7Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B764));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R0_INV_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y7__R1_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B50));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R1_INV_0 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R2_INV_0 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R2_INV_1 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B836));
  sky130_fd_sc_hd__clkbuf_4 T7Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8647));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R0_INV_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8683));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R1_INV_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R2_INV_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R2_INV_1 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y80__R3_BUF_0 (.A(clk_L1_B544), .X(clk_L0_B8719));
  sky130_fd_sc_hd__clkbuf_4 T7Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8755));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R0_INV_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8791));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R1_INV_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R2_INV_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R2_INV_1 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8827));
  sky130_fd_sc_hd__clkbuf_4 T7Y82__R0_BUF_0 (.A(clk_L1_B553), .X(clk_L0_B8863));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R0_INV_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8899));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R1_INV_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R2_INV_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R2_INV_1 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8935));
  sky130_fd_sc_hd__clkbuf_4 T7Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8971));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R0_INV_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y83__R1_BUF_0 (.A(clk_L1_B562), .X(clk_L0_B9007));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R1_INV_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R2_INV_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R2_INV_1 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9043));
  sky130_fd_sc_hd__clkbuf_4 T7Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9079));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R0_INV_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9115));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R1_INV_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R2_INV_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R2_INV_1 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y84__R3_BUF_0 (.A(clk_L1_B571), .X(clk_L0_B9151));
  sky130_fd_sc_hd__clkbuf_4 T7Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9187));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R0_INV_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9223));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R1_INV_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R2_INV_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R2_INV_1 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9259));
  sky130_fd_sc_hd__clkbuf_4 T7Y86__R0_BUF_0 (.A(clk_L1_B580), .X(clk_L0_B9295));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R0_INV_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9331));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R1_INV_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R2_INV_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R2_INV_1 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9367));
  sky130_fd_sc_hd__clkbuf_4 T7Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9403));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R0_INV_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y87__R1_BUF_0 (.A(clk_L1_B589), .X(clk_L0_B9439));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R1_INV_0 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R2_INV_0 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R2_INV_1 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9475));
  sky130_fd_sc_hd__clkbuf_4 T7Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9511));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R0_INV_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9547));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R1_INV_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R2_INV_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R2_INV_1 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y88__R3_BUF_0 (.A(clk_L1_B598), .X(clk_L0_B9583));
  sky130_fd_sc_hd__clkbuf_4 T7Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9619));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R0_INV_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9655));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R1_INV_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R2_INV_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R2_INV_1 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9691));
  sky130_fd_sc_hd__clkbuf_4 T7Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B872));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R0_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B908));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R1_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R2_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R2_INV_1 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y8__R3_BUF_0 (.A(clk_L2_B3), .X(clk_L1_B59));
  sky130_fd_sc_hd__clkbuf_4 T7Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B980));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R0_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1016));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R1_INV_0 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R2_INV_0 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R2_INV_1 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1052));
  sky130_fd_sc_hd__clkbuf_4 T8Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B18));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R0_INV_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B53));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R1_INV_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R2_INV_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R2_INV_1 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B88));
  sky130_fd_sc_hd__clkbuf_4 T8Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1089));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R0_INV_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1125));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R1_INV_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R2_INV_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R2_INV_1 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1161));
  sky130_fd_sc_hd__clkbuf_4 T8Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1197));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R0_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1233));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R1_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R2_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R2_INV_1 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1269));
  sky130_fd_sc_hd__clkbuf_4 T8Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1305));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R0_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1341));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R1_INV_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R2_INV_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R2_INV_1 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1377));
  sky130_fd_sc_hd__clkbuf_4 T8Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1413));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R0_INV_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1449));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R1_INV_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R2_INV_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R2_INV_1 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1485));
  sky130_fd_sc_hd__clkbuf_4 T8Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1521));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R0_INV_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1556));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R1_INV_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R2_INV_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R2_INV_1 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1592));
  sky130_fd_sc_hd__clkbuf_4 T8Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1628));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R0_INV_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y15__R1_BUF_0 (.A(clk_L2_B6), .X(clk_L1_B104));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R1_INV_0 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R2_INV_0 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R2_INV_1 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1700));
  sky130_fd_sc_hd__clkbuf_4 T8Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1736));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R0_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1772));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R1_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R2_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R2_INV_1 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y16__R3_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B113));
  sky130_fd_sc_hd__clkbuf_4 T8Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1844));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R0_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1880));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R1_INV_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R2_INV_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R2_INV_1 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1916));
  sky130_fd_sc_hd__clkbuf_4 T8Y18__R0_BUF_0 (.A(clk_L2_B7), .X(clk_L1_B122));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R0_INV_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1988));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R1_INV_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R2_INV_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R2_INV_1 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2024));
  sky130_fd_sc_hd__clkbuf_4 T8Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2060));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R0_INV_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y19__R1_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B131));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R1_INV_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R2_INV_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R2_INV_1 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2132));
  sky130_fd_sc_hd__clkbuf_4 T8Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B123));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R0_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B158));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R1_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R2_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R2_INV_1 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B193));
  sky130_fd_sc_hd__clkbuf_4 T8Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2168));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R0_INV_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2204));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R1_INV_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R2_INV_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R2_INV_1 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y20__R3_BUF_0 (.A(clk_L2_B8), .X(clk_L1_B140));
  sky130_fd_sc_hd__clkbuf_4 T8Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2276));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R0_INV_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2312));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R1_INV_0 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R2_INV_0 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R2_INV_1 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2348));
  sky130_fd_sc_hd__clkbuf_4 T8Y22__R0_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B149));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R0_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2420));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R1_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R2_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R2_INV_1 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2456));
  sky130_fd_sc_hd__clkbuf_4 T8Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2492));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R0_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y23__R1_BUF_0 (.A(clk_L2_B9), .X(clk_L1_B158));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R1_INV_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R2_INV_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R2_INV_1 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2564));
  sky130_fd_sc_hd__clkbuf_4 T8Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2600));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R0_INV_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2636));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R1_INV_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R2_INV_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R2_INV_1 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y24__R3_BUF_0 (.A(clk_L2_B10), .X(clk_L1_B167));
  sky130_fd_sc_hd__clkbuf_4 T8Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2708));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R0_INV_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2744));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R1_INV_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R2_INV_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R2_INV_1 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2780));
  sky130_fd_sc_hd__clkbuf_4 T8Y26__R0_BUF_0 (.A(clk_L3_B0), .X(clk_L2_B11));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R0_INV_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2852));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R1_INV_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R2_INV_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R2_INV_1 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2888));
  sky130_fd_sc_hd__clkbuf_4 T8Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2924));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R0_INV_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y27__R1_BUF_0 (.A(clk_L2_B11), .X(clk_L1_B185));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R1_INV_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R2_INV_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R2_INV_1 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2996));
  sky130_fd_sc_hd__clkbuf_4 T8Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3032));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R0_INV_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3068));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R1_INV_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R2_INV_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R2_INV_1 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y28__R3_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B194));
  sky130_fd_sc_hd__clkbuf_4 T8Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3140));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R0_INV_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3176));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R1_INV_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R2_INV_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R2_INV_1 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3212));
  sky130_fd_sc_hd__clkbuf_4 T8Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B228));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R0_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B263));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R1_INV_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R2_INV_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R2_INV_1 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B299));
  sky130_fd_sc_hd__clkbuf_4 T8Y30__R0_BUF_0 (.A(clk_L2_B12), .X(clk_L1_B203));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R0_INV_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3284));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R1_INV_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R2_INV_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R2_INV_1 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3320));
  sky130_fd_sc_hd__clkbuf_4 T8Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3356));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R0_INV_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y31__R1_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B212));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R1_INV_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R2_INV_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R2_INV_1 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3428));
  sky130_fd_sc_hd__clkbuf_4 T8Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3464));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R0_INV_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3500));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R1_INV_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R2_INV_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R2_INV_1 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y32__R3_BUF_0 (.A(clk_L2_B13), .X(clk_L1_B221));
  sky130_fd_sc_hd__clkbuf_4 T8Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3572));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R0_INV_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3608));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R1_INV_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R2_INV_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R2_INV_1 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3644));
  sky130_fd_sc_hd__clkbuf_4 T8Y34__R0_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B230));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R0_INV_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3716));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R1_INV_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R2_INV_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R2_INV_1 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3752));
  sky130_fd_sc_hd__clkbuf_4 T8Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3788));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R0_INV_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y35__R1_BUF_0 (.A(clk_L2_B14), .X(clk_L1_B239));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R1_INV_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R2_INV_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R2_INV_1 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3860));
  sky130_fd_sc_hd__clkbuf_4 T8Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3896));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R0_INV_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3932));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R1_INV_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R2_INV_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R2_INV_1 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y36__R3_BUF_0 (.A(clk_L2_B15), .X(clk_L1_B248));
  sky130_fd_sc_hd__clkbuf_4 T8Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4004));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R0_INV_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4040));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R1_INV_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R2_INV_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R2_INV_1 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4076));
  sky130_fd_sc_hd__clkbuf_4 T8Y38__R0_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B257));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R0_INV_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4148));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R1_INV_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R2_INV_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R2_INV_1 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4184));
  sky130_fd_sc_hd__clkbuf_4 T8Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4220));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R0_INV_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y39__R1_BUF_0 (.A(clk_L2_B16), .X(clk_L1_B266));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R1_INV_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R2_INV_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R2_INV_1 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4292));
  sky130_fd_sc_hd__clkbuf_4 T8Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B334));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R0_INV_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B369));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R1_INV_0 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R2_INV_0 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R2_INV_1 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B405));
  sky130_fd_sc_hd__clkbuf_4 T8Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4328));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R0_INV_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4364));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R1_INV_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R2_INV_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R2_INV_1 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y40__R3_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B275));
  sky130_fd_sc_hd__clkbuf_4 T8Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4436));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R0_INV_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4472));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R1_INV_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R2_INV_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R2_INV_1 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4508));
  sky130_fd_sc_hd__clkbuf_4 T8Y42__R0_BUF_0 (.A(clk_L2_B17), .X(clk_L1_B284));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R0_INV_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4580));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R1_INV_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R2_INV_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R2_INV_1 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4616));
  sky130_fd_sc_hd__clkbuf_4 T8Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4652));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R0_INV_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y43__R1_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B293));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R1_INV_0 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R2_INV_0 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R2_INV_1 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4724));
  sky130_fd_sc_hd__clkbuf_4 T8Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4760));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R0_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4796));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R1_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R2_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R2_INV_1 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y44__R3_BUF_0 (.A(clk_L2_B18), .X(clk_L1_B302));
  sky130_fd_sc_hd__clkbuf_4 T8Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4868));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R0_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4904));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R1_INV_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R2_INV_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R2_INV_1 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4940));
  sky130_fd_sc_hd__clkbuf_4 T8Y46__R0_BUF_0 (.A(clk_L2_B19), .X(clk_L1_B311));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R0_INV_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5012));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R1_INV_0 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R2_INV_0 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R2_INV_1 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5048));
  sky130_fd_sc_hd__clkbuf_4 T8Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5084));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R0_INV_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y47__R1_BUF_0 (.A(clk_L3_B1), .X(clk_L2_B20));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R1_INV_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R2_INV_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R2_INV_1 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5156));
  sky130_fd_sc_hd__clkbuf_4 T8Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5192));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R0_INV_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5228));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R1_INV_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R2_INV_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R2_INV_1 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y48__R3_BUF_0 (.A(clk_L2_B20), .X(clk_L1_B329));
  sky130_fd_sc_hd__clkbuf_4 T8Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5300));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R0_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5336));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R1_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R2_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R2_INV_1 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5372));
  sky130_fd_sc_hd__clkbuf_4 T8Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B441));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R0_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B477));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R1_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R2_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R2_INV_1 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B513));
  sky130_fd_sc_hd__clkbuf_4 T8Y50__R0_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B338));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R0_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5444));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R1_INV_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R2_INV_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R2_INV_1 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5480));
  sky130_fd_sc_hd__clkbuf_4 T8Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5516));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R0_INV_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y51__R1_BUF_0 (.A(clk_L2_B21), .X(clk_L1_B347));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R1_INV_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R2_INV_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R2_INV_1 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5588));
  sky130_fd_sc_hd__clkbuf_4 T8Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5624));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R0_INV_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5660));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R1_INV_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R2_INV_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R2_INV_1 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y52__R3_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B356));
  sky130_fd_sc_hd__clkbuf_4 T8Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5732));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R0_INV_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5768));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R1_INV_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R2_INV_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R2_INV_1 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5804));
  sky130_fd_sc_hd__clkbuf_4 T8Y54__R0_BUF_0 (.A(clk_L2_B22), .X(clk_L1_B365));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R0_INV_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5876));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R1_INV_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R2_INV_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R2_INV_1 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5912));
  sky130_fd_sc_hd__clkbuf_4 T8Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5948));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R0_INV_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y55__R1_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B374));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R1_INV_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R2_INV_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R2_INV_1 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6020));
  sky130_fd_sc_hd__clkbuf_4 T8Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6056));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R0_INV_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6092));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R1_INV_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R2_INV_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R2_INV_1 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y56__R3_BUF_0 (.A(clk_L2_B23), .X(clk_L1_B383));
  sky130_fd_sc_hd__clkbuf_4 T8Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6164));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R0_INV_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6200));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R1_INV_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R2_INV_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R2_INV_1 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6236));
  sky130_fd_sc_hd__clkbuf_4 T8Y58__R0_BUF_0 (.A(clk_L2_B24), .X(clk_L1_B392));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R0_INV_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6308));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R1_INV_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R2_INV_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R2_INV_1 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6344));
  sky130_fd_sc_hd__clkbuf_4 T8Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6380));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R0_INV_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y59__R1_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B401));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R1_INV_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R2_INV_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R2_INV_1 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6452));
  sky130_fd_sc_hd__clkbuf_4 T8Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B549));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R0_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B585));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R1_INV_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R2_INV_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R2_INV_1 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B621));
  sky130_fd_sc_hd__clkbuf_4 T8Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6488));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R0_INV_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6524));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R1_INV_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R2_INV_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R2_INV_1 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y60__R3_BUF_0 (.A(clk_L2_B25), .X(clk_L1_B410));
  sky130_fd_sc_hd__clkbuf_4 T8Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6596));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R0_INV_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6632));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R1_INV_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R2_INV_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R2_INV_1 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6668));
  sky130_fd_sc_hd__clkbuf_4 T8Y62__R0_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B419));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R0_INV_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6740));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R1_INV_0 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R2_INV_0 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R2_INV_1 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6776));
  sky130_fd_sc_hd__clkbuf_4 T8Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6812));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R0_INV_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y63__R1_BUF_0 (.A(clk_L2_B26), .X(clk_L1_B428));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R1_INV_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R2_INV_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R2_INV_1 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6884));
  sky130_fd_sc_hd__clkbuf_4 T8Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6920));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R0_INV_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6956));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R1_INV_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R2_INV_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R2_INV_1 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y64__R3_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B437));
  sky130_fd_sc_hd__clkbuf_4 T8Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7028));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R0_INV_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7064));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R1_INV_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R2_INV_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R2_INV_1 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7100));
  sky130_fd_sc_hd__clkbuf_4 T8Y66__R0_BUF_0 (.A(clk_L2_B27), .X(clk_L1_B446));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R0_INV_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7172));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R1_INV_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R2_INV_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R2_INV_1 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7208));
  sky130_fd_sc_hd__clkbuf_4 T8Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7244));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R0_INV_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y67__R1_BUF_0 (.A(clk_L2_B28), .X(clk_L1_B455));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R1_INV_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R2_INV_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R2_INV_1 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7316));
  sky130_fd_sc_hd__clkbuf_4 T8Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7352));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R0_INV_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7388));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R1_INV_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R2_INV_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R2_INV_1 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y68__R3_BUF_0 (.A(clk_L3_B2), .X(clk_L2_B29));
  sky130_fd_sc_hd__clkbuf_4 T8Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7460));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R0_INV_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7496));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R1_INV_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R2_INV_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R2_INV_1 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7532));
  sky130_fd_sc_hd__clkbuf_4 T8Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B657));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R0_INV_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B693));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R1_INV_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R2_INV_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R2_INV_1 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B729));
  sky130_fd_sc_hd__clkbuf_4 T8Y70__R0_BUF_0 (.A(clk_L2_B29), .X(clk_L1_B473));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R0_INV_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7604));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R1_INV_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R2_INV_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R2_INV_1 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7640));
  sky130_fd_sc_hd__clkbuf_4 T8Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7676));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R0_INV_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y71__R1_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B482));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R1_INV_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R2_INV_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R2_INV_1 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7748));
  sky130_fd_sc_hd__clkbuf_4 T8Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7784));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R0_INV_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7820));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R1_INV_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R2_INV_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R2_INV_1 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y72__R3_BUF_0 (.A(clk_L2_B30), .X(clk_L1_B491));
  sky130_fd_sc_hd__clkbuf_4 T8Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7892));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R0_INV_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7928));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R1_INV_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R2_INV_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R2_INV_1 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7964));
  sky130_fd_sc_hd__clkbuf_4 T8Y74__R0_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B500));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R0_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8036));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R1_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R2_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R2_INV_1 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8072));
  sky130_fd_sc_hd__clkbuf_4 T8Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8108));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R0_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y75__R1_BUF_0 (.A(clk_L2_B31), .X(clk_L1_B509));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R1_INV_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R2_INV_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R2_INV_1 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8180));
  sky130_fd_sc_hd__clkbuf_4 T8Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8216));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R0_INV_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8252));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R1_INV_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R2_INV_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R2_INV_1 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y76__R3_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B518));
  sky130_fd_sc_hd__clkbuf_4 T8Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8324));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R0_INV_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8360));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R1_INV_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R2_INV_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R2_INV_1 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8396));
  sky130_fd_sc_hd__clkbuf_4 T8Y78__R0_BUF_0 (.A(clk_L2_B32), .X(clk_L1_B527));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R0_INV_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8468));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R1_INV_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R2_INV_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R2_INV_1 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8504));
  sky130_fd_sc_hd__clkbuf_4 T8Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8540));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R0_INV_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y79__R1_BUF_0 (.A(clk_L2_B33), .X(clk_L1_B536));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R1_INV_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R2_INV_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R2_INV_1 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8612));
  sky130_fd_sc_hd__clkbuf_4 T8Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B765));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R0_INV_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B801));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R1_INV_0 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R2_INV_0 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R2_INV_1 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B837));
  sky130_fd_sc_hd__clkbuf_4 T8Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8648));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R0_INV_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8684));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R1_INV_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R2_INV_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R2_INV_1 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y80__R3_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B545));
  sky130_fd_sc_hd__clkbuf_4 T8Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8756));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R0_INV_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8792));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R1_INV_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R2_INV_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R2_INV_1 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8828));
  sky130_fd_sc_hd__clkbuf_4 T8Y82__R0_BUF_0 (.A(clk_L2_B34), .X(clk_L1_B554));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R0_INV_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8900));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R1_INV_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R2_INV_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R2_INV_1 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8936));
  sky130_fd_sc_hd__clkbuf_4 T8Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8972));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R0_INV_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y83__R1_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B563));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R1_INV_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R2_INV_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R2_INV_1 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9044));
  sky130_fd_sc_hd__clkbuf_4 T8Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9080));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R0_INV_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9116));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R1_INV_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R2_INV_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R2_INV_1 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y84__R3_BUF_0 (.A(clk_L2_B35), .X(clk_L1_B572));
  sky130_fd_sc_hd__clkbuf_4 T8Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9188));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R0_INV_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9224));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R1_INV_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R2_INV_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R2_INV_1 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9260));
  sky130_fd_sc_hd__clkbuf_4 T8Y86__R0_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B581));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R0_INV_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9332));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R1_INV_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R2_INV_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R2_INV_1 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9368));
  sky130_fd_sc_hd__clkbuf_4 T8Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9404));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R0_INV_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y87__R1_BUF_0 (.A(clk_L2_B36), .X(clk_L1_B590));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R1_INV_0 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R2_INV_0 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R2_INV_1 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9476));
  sky130_fd_sc_hd__clkbuf_4 T8Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9512));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R0_INV_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9548));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R1_INV_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R2_INV_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R2_INV_1 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y88__R3_BUF_0 (.A(clk_L2_B37), .X(clk_L1_B599));
  sky130_fd_sc_hd__clkbuf_4 T8Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9620));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R0_INV_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9656));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R1_INV_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R2_INV_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R2_INV_1 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9692));
  sky130_fd_sc_hd__clkbuf_4 T8Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B873));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R0_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B909));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R1_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R2_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R2_INV_1 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B945));
  sky130_fd_sc_hd__clkbuf_4 T8Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B981));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R0_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1017));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R1_INV_0 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R2_INV_0 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R2_INV_1 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1053));
  sky130_fd_sc_hd__clkbuf_4 T9Y0__R0_BUF_0 (.A(clk_L1_B1), .X(clk_L0_B19));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R0_INV_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y0__R1_BUF_0 (.A(clk_L1_B3), .X(clk_L0_B54));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R1_INV_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R2_INV_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R2_INV_1 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y0__R3_BUF_0 (.A(clk_L1_B5), .X(clk_L0_B89));
  sky130_fd_sc_hd__clkbuf_4 T9Y10__R0_BUF_0 (.A(clk_L1_B68), .X(clk_L0_B1090));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R0_INV_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y10__R1_BUF_0 (.A(clk_L1_B70), .X(clk_L0_B1126));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R1_INV_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R2_INV_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R2_INV_1 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y10__R3_BUF_0 (.A(clk_L1_B72), .X(clk_L0_B1162));
  sky130_fd_sc_hd__clkbuf_4 T9Y11__R0_BUF_0 (.A(clk_L1_B74), .X(clk_L0_B1198));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R0_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y11__R1_BUF_0 (.A(clk_L1_B77), .X(clk_L0_B1234));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R1_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R2_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R2_INV_1 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y11__R3_BUF_0 (.A(clk_L1_B79), .X(clk_L0_B1270));
  sky130_fd_sc_hd__clkbuf_4 T9Y12__R0_BUF_0 (.A(clk_L1_B81), .X(clk_L0_B1306));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R0_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y12__R1_BUF_0 (.A(clk_L1_B83), .X(clk_L0_B1342));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R1_INV_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R2_INV_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R2_INV_1 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y12__R3_BUF_0 (.A(clk_L1_B86), .X(clk_L0_B1378));
  sky130_fd_sc_hd__clkbuf_4 T9Y13__R0_BUF_0 (.A(clk_L1_B88), .X(clk_L0_B1414));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R0_INV_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y13__R1_BUF_0 (.A(clk_L1_B90), .X(clk_L0_B1450));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R1_INV_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R2_INV_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R2_INV_1 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y13__R3_BUF_0 (.A(clk_L1_B92), .X(clk_L0_B1486));
  sky130_fd_sc_hd__clkbuf_4 T9Y14__R0_BUF_0 (.A(clk_L1_B95), .X(clk_L0_B1522));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R0_INV_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y14__R1_BUF_0 (.A(clk_L1_B97), .X(clk_L0_B1557));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R1_INV_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R2_INV_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R2_INV_1 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y14__R3_BUF_0 (.A(clk_L1_B99), .X(clk_L0_B1593));
  sky130_fd_sc_hd__clkbuf_4 T9Y15__R0_BUF_0 (.A(clk_L1_B101), .X(clk_L0_B1629));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R0_INV_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y15__R1_BUF_0 (.A(clk_L1_B104), .X(clk_L0_B1665));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R1_INV_0 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R2_INV_0 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R2_INV_1 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y15__R3_BUF_0 (.A(clk_L1_B106), .X(clk_L0_B1701));
  sky130_fd_sc_hd__clkbuf_4 T9Y16__R0_BUF_0 (.A(clk_L1_B108), .X(clk_L0_B1737));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R0_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y16__R1_BUF_0 (.A(clk_L1_B110), .X(clk_L0_B1773));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R1_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R2_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R2_INV_1 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y16__R3_BUF_0 (.A(clk_L1_B113), .X(clk_L0_B1809));
  sky130_fd_sc_hd__clkbuf_4 T9Y17__R0_BUF_0 (.A(clk_L1_B115), .X(clk_L0_B1845));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R0_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y17__R1_BUF_0 (.A(clk_L1_B117), .X(clk_L0_B1881));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R1_INV_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R2_INV_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R2_INV_1 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y17__R3_BUF_0 (.A(clk_L1_B119), .X(clk_L0_B1917));
  sky130_fd_sc_hd__clkbuf_4 T9Y18__R0_BUF_0 (.A(clk_L1_B122), .X(clk_L0_B1953));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R0_INV_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y18__R1_BUF_0 (.A(clk_L1_B124), .X(clk_L0_B1989));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R1_INV_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R2_INV_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R2_INV_1 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y18__R3_BUF_0 (.A(clk_L1_B126), .X(clk_L0_B2025));
  sky130_fd_sc_hd__clkbuf_4 T9Y19__R0_BUF_0 (.A(clk_L1_B128), .X(clk_L0_B2061));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R0_INV_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y19__R1_BUF_0 (.A(clk_L1_B131), .X(clk_L0_B2097));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R1_INV_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R2_INV_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R2_INV_1 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y19__R3_BUF_0 (.A(clk_L1_B133), .X(clk_L0_B2133));
  sky130_fd_sc_hd__clkbuf_4 T9Y1__R0_BUF_0 (.A(clk_L1_B7), .X(clk_L0_B124));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R0_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y1__R1_BUF_0 (.A(clk_L1_B9), .X(clk_L0_B159));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R1_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R2_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R2_INV_1 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y1__R3_BUF_0 (.A(clk_L1_B12), .X(clk_L0_B194));
  sky130_fd_sc_hd__clkbuf_4 T9Y20__R0_BUF_0 (.A(clk_L1_B135), .X(clk_L0_B2169));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R0_INV_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y20__R1_BUF_0 (.A(clk_L1_B137), .X(clk_L0_B2205));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R1_INV_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R2_INV_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R2_INV_1 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y20__R3_BUF_0 (.A(clk_L1_B140), .X(clk_L0_B2241));
  sky130_fd_sc_hd__clkbuf_4 T9Y21__R0_BUF_0 (.A(clk_L1_B142), .X(clk_L0_B2277));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R0_INV_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y21__R1_BUF_0 (.A(clk_L1_B144), .X(clk_L0_B2313));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R1_INV_0 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R2_INV_0 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R2_INV_1 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y21__R3_BUF_0 (.A(clk_L1_B146), .X(clk_L0_B2349));
  sky130_fd_sc_hd__clkbuf_4 T9Y22__R0_BUF_0 (.A(clk_L1_B149), .X(clk_L0_B2385));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R0_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y22__R1_BUF_0 (.A(clk_L1_B151), .X(clk_L0_B2421));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R1_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R2_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R2_INV_1 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y22__R3_BUF_0 (.A(clk_L1_B153), .X(clk_L0_B2457));
  sky130_fd_sc_hd__clkbuf_4 T9Y23__R0_BUF_0 (.A(clk_L1_B155), .X(clk_L0_B2493));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R0_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y23__R1_BUF_0 (.A(clk_L1_B158), .X(clk_L0_B2529));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R1_INV_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R2_INV_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R2_INV_1 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y23__R3_BUF_0 (.A(clk_L1_B160), .X(clk_L0_B2565));
  sky130_fd_sc_hd__clkbuf_4 T9Y24__R0_BUF_0 (.A(clk_L1_B162), .X(clk_L0_B2601));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R0_INV_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y24__R1_BUF_0 (.A(clk_L1_B164), .X(clk_L0_B2637));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R1_INV_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R2_INV_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R2_INV_1 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y24__R3_BUF_0 (.A(clk_L1_B167), .X(clk_L0_B2673));
  sky130_fd_sc_hd__clkbuf_4 T9Y25__R0_BUF_0 (.A(clk_L1_B169), .X(clk_L0_B2709));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R0_INV_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y25__R1_BUF_0 (.A(clk_L1_B171), .X(clk_L0_B2745));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R1_INV_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R2_INV_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R2_INV_1 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y25__R3_BUF_0 (.A(clk_L1_B173), .X(clk_L0_B2781));
  sky130_fd_sc_hd__clkbuf_4 T9Y26__R0_BUF_0 (.A(clk_L1_B176), .X(clk_L0_B2817));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R0_INV_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y26__R1_BUF_0 (.A(clk_L1_B178), .X(clk_L0_B2853));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R1_INV_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R2_INV_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R2_INV_1 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y26__R3_BUF_0 (.A(clk_L1_B180), .X(clk_L0_B2889));
  sky130_fd_sc_hd__clkbuf_4 T9Y27__R0_BUF_0 (.A(clk_L1_B182), .X(clk_L0_B2925));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R0_INV_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y27__R1_BUF_0 (.A(clk_L1_B185), .X(clk_L0_B2961));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R1_INV_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R2_INV_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R2_INV_1 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y27__R3_BUF_0 (.A(clk_L1_B187), .X(clk_L0_B2997));
  sky130_fd_sc_hd__clkbuf_4 T9Y28__R0_BUF_0 (.A(clk_L1_B189), .X(clk_L0_B3033));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R0_INV_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y28__R1_BUF_0 (.A(clk_L1_B191), .X(clk_L0_B3069));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R1_INV_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R2_INV_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R2_INV_1 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y28__R3_BUF_0 (.A(clk_L1_B194), .X(clk_L0_B3105));
  sky130_fd_sc_hd__clkbuf_4 T9Y29__R0_BUF_0 (.A(clk_L1_B196), .X(clk_L0_B3141));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R0_INV_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y29__R1_BUF_0 (.A(clk_L1_B198), .X(clk_L0_B3177));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R1_INV_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R2_INV_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R2_INV_1 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y29__R3_BUF_0 (.A(clk_L1_B200), .X(clk_L0_B3213));
  sky130_fd_sc_hd__clkbuf_4 T9Y2__R0_BUF_0 (.A(clk_L1_B14), .X(clk_L0_B229));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R0_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y2__R1_BUF_0 (.A(clk_L1_B16), .X(clk_L0_B264));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R1_INV_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R2_INV_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R2_INV_1 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y2__R3_BUF_0 (.A(clk_L1_B18), .X(clk_L0_B300));
  sky130_fd_sc_hd__clkbuf_4 T9Y30__R0_BUF_0 (.A(clk_L1_B203), .X(clk_L0_B3249));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R0_INV_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y30__R1_BUF_0 (.A(clk_L1_B205), .X(clk_L0_B3285));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R1_INV_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R2_INV_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R2_INV_1 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y30__R3_BUF_0 (.A(clk_L1_B207), .X(clk_L0_B3321));
  sky130_fd_sc_hd__clkbuf_4 T9Y31__R0_BUF_0 (.A(clk_L1_B209), .X(clk_L0_B3357));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R0_INV_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y31__R1_BUF_0 (.A(clk_L1_B212), .X(clk_L0_B3393));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R1_INV_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R2_INV_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R2_INV_1 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y31__R3_BUF_0 (.A(clk_L1_B214), .X(clk_L0_B3429));
  sky130_fd_sc_hd__clkbuf_4 T9Y32__R0_BUF_0 (.A(clk_L1_B216), .X(clk_L0_B3465));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R0_INV_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y32__R1_BUF_0 (.A(clk_L1_B218), .X(clk_L0_B3501));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R1_INV_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R2_INV_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R2_INV_1 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y32__R3_BUF_0 (.A(clk_L1_B221), .X(clk_L0_B3537));
  sky130_fd_sc_hd__clkbuf_4 T9Y33__R0_BUF_0 (.A(clk_L1_B223), .X(clk_L0_B3573));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R0_INV_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y33__R1_BUF_0 (.A(clk_L1_B225), .X(clk_L0_B3609));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R1_INV_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R2_INV_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R2_INV_1 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y33__R3_BUF_0 (.A(clk_L1_B227), .X(clk_L0_B3645));
  sky130_fd_sc_hd__clkbuf_4 T9Y34__R0_BUF_0 (.A(clk_L1_B230), .X(clk_L0_B3681));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R0_INV_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y34__R1_BUF_0 (.A(clk_L1_B232), .X(clk_L0_B3717));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R1_INV_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R2_INV_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R2_INV_1 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y34__R3_BUF_0 (.A(clk_L1_B234), .X(clk_L0_B3753));
  sky130_fd_sc_hd__clkbuf_4 T9Y35__R0_BUF_0 (.A(clk_L1_B236), .X(clk_L0_B3789));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R0_INV_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y35__R1_BUF_0 (.A(clk_L1_B239), .X(clk_L0_B3825));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R1_INV_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R2_INV_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R2_INV_1 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y35__R3_BUF_0 (.A(clk_L1_B241), .X(clk_L0_B3861));
  sky130_fd_sc_hd__clkbuf_4 T9Y36__R0_BUF_0 (.A(clk_L1_B243), .X(clk_L0_B3897));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R0_INV_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y36__R1_BUF_0 (.A(clk_L1_B245), .X(clk_L0_B3933));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R1_INV_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R2_INV_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R2_INV_1 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y36__R3_BUF_0 (.A(clk_L1_B248), .X(clk_L0_B3969));
  sky130_fd_sc_hd__clkbuf_4 T9Y37__R0_BUF_0 (.A(clk_L1_B250), .X(clk_L0_B4005));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R0_INV_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y37__R1_BUF_0 (.A(clk_L1_B252), .X(clk_L0_B4041));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R1_INV_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R2_INV_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R2_INV_1 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y37__R3_BUF_0 (.A(clk_L1_B254), .X(clk_L0_B4077));
  sky130_fd_sc_hd__clkbuf_4 T9Y38__R0_BUF_0 (.A(clk_L1_B257), .X(clk_L0_B4113));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R0_INV_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y38__R1_BUF_0 (.A(clk_L1_B259), .X(clk_L0_B4149));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R1_INV_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R2_INV_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R2_INV_1 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y38__R3_BUF_0 (.A(clk_L1_B261), .X(clk_L0_B4185));
  sky130_fd_sc_hd__clkbuf_4 T9Y39__R0_BUF_0 (.A(clk_L1_B263), .X(clk_L0_B4221));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R0_INV_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y39__R1_BUF_0 (.A(clk_L1_B266), .X(clk_L0_B4257));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R1_INV_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R2_INV_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R2_INV_1 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y39__R3_BUF_0 (.A(clk_L1_B268), .X(clk_L0_B4293));
  sky130_fd_sc_hd__clkbuf_4 T9Y3__R0_BUF_0 (.A(clk_L1_B20), .X(clk_L0_B335));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R0_INV_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y3__R1_BUF_0 (.A(clk_L1_B23), .X(clk_L0_B370));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R1_INV_0 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R2_INV_0 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R2_INV_1 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y3__R3_BUF_0 (.A(clk_L1_B25), .X(clk_L0_B406));
  sky130_fd_sc_hd__clkbuf_4 T9Y40__R0_BUF_0 (.A(clk_L1_B270), .X(clk_L0_B4329));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R0_INV_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y40__R1_BUF_0 (.A(clk_L1_B272), .X(clk_L0_B4365));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R1_INV_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R2_INV_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R2_INV_1 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y40__R3_BUF_0 (.A(clk_L1_B275), .X(clk_L0_B4401));
  sky130_fd_sc_hd__clkbuf_4 T9Y41__R0_BUF_0 (.A(clk_L1_B277), .X(clk_L0_B4437));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R0_INV_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y41__R1_BUF_0 (.A(clk_L1_B279), .X(clk_L0_B4473));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R1_INV_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R2_INV_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R2_INV_1 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y41__R3_BUF_0 (.A(clk_L1_B281), .X(clk_L0_B4509));
  sky130_fd_sc_hd__clkbuf_4 T9Y42__R0_BUF_0 (.A(clk_L1_B284), .X(clk_L0_B4545));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R0_INV_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y42__R1_BUF_0 (.A(clk_L1_B286), .X(clk_L0_B4581));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R1_INV_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R2_INV_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R2_INV_1 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y42__R3_BUF_0 (.A(clk_L1_B288), .X(clk_L0_B4617));
  sky130_fd_sc_hd__clkbuf_4 T9Y43__R0_BUF_0 (.A(clk_L1_B290), .X(clk_L0_B4653));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R0_INV_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y43__R1_BUF_0 (.A(clk_L1_B293), .X(clk_L0_B4689));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R1_INV_0 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R2_INV_0 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R2_INV_1 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y43__R3_BUF_0 (.A(clk_L1_B295), .X(clk_L0_B4725));
  sky130_fd_sc_hd__clkbuf_4 T9Y44__R0_BUF_0 (.A(clk_L1_B297), .X(clk_L0_B4761));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R0_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y44__R1_BUF_0 (.A(clk_L1_B299), .X(clk_L0_B4797));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R1_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R2_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R2_INV_1 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y44__R3_BUF_0 (.A(clk_L1_B302), .X(clk_L0_B4833));
  sky130_fd_sc_hd__clkbuf_4 T9Y45__R0_BUF_0 (.A(clk_L1_B304), .X(clk_L0_B4869));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R0_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y45__R1_BUF_0 (.A(clk_L1_B306), .X(clk_L0_B4905));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R1_INV_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R2_INV_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R2_INV_1 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y45__R3_BUF_0 (.A(clk_L1_B308), .X(clk_L0_B4941));
  sky130_fd_sc_hd__clkbuf_4 T9Y46__R0_BUF_0 (.A(clk_L1_B311), .X(clk_L0_B4977));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R0_INV_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y46__R1_BUF_0 (.A(clk_L1_B313), .X(clk_L0_B5013));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R1_INV_0 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R2_INV_0 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R2_INV_1 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y46__R3_BUF_0 (.A(clk_L1_B315), .X(clk_L0_B5049));
  sky130_fd_sc_hd__clkbuf_4 T9Y47__R0_BUF_0 (.A(clk_L1_B317), .X(clk_L0_B5085));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R0_INV_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y47__R1_BUF_0 (.A(clk_L1_B320), .X(clk_L0_B5121));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R1_INV_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R2_INV_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R2_INV_1 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y47__R3_BUF_0 (.A(clk_L1_B322), .X(clk_L0_B5157));
  sky130_fd_sc_hd__clkbuf_4 T9Y48__R0_BUF_0 (.A(clk_L1_B324), .X(clk_L0_B5193));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R0_INV_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y48__R1_BUF_0 (.A(clk_L1_B326), .X(clk_L0_B5229));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R1_INV_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R2_INV_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R2_INV_1 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y48__R3_BUF_0 (.A(clk_L1_B329), .X(clk_L0_B5265));
  sky130_fd_sc_hd__clkbuf_4 T9Y49__R0_BUF_0 (.A(clk_L1_B331), .X(clk_L0_B5301));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R0_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y49__R1_BUF_0 (.A(clk_L1_B333), .X(clk_L0_B5337));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R1_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R2_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R2_INV_1 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y49__R3_BUF_0 (.A(clk_L1_B335), .X(clk_L0_B5373));
  sky130_fd_sc_hd__clkbuf_4 T9Y4__R0_BUF_0 (.A(clk_L1_B27), .X(clk_L0_B442));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R0_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y4__R1_BUF_0 (.A(clk_L1_B29), .X(clk_L0_B478));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R1_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R2_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R2_INV_1 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y4__R3_BUF_0 (.A(clk_L1_B32), .X(clk_L0_B514));
  sky130_fd_sc_hd__clkbuf_4 T9Y50__R0_BUF_0 (.A(clk_L1_B338), .X(clk_L0_B5409));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R0_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y50__R1_BUF_0 (.A(clk_L1_B340), .X(clk_L0_B5445));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R1_INV_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R2_INV_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R2_INV_1 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y50__R3_BUF_0 (.A(clk_L1_B342), .X(clk_L0_B5481));
  sky130_fd_sc_hd__clkbuf_4 T9Y51__R0_BUF_0 (.A(clk_L1_B344), .X(clk_L0_B5517));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R0_INV_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y51__R1_BUF_0 (.A(clk_L1_B347), .X(clk_L0_B5553));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R1_INV_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R2_INV_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R2_INV_1 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y51__R3_BUF_0 (.A(clk_L1_B349), .X(clk_L0_B5589));
  sky130_fd_sc_hd__clkbuf_4 T9Y52__R0_BUF_0 (.A(clk_L1_B351), .X(clk_L0_B5625));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R0_INV_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y52__R1_BUF_0 (.A(clk_L1_B353), .X(clk_L0_B5661));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R1_INV_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R2_INV_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R2_INV_1 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y52__R3_BUF_0 (.A(clk_L1_B356), .X(clk_L0_B5697));
  sky130_fd_sc_hd__clkbuf_4 T9Y53__R0_BUF_0 (.A(clk_L1_B358), .X(clk_L0_B5733));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R0_INV_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y53__R1_BUF_0 (.A(clk_L1_B360), .X(clk_L0_B5769));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R1_INV_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R2_INV_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R2_INV_1 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y53__R3_BUF_0 (.A(clk_L1_B362), .X(clk_L0_B5805));
  sky130_fd_sc_hd__clkbuf_4 T9Y54__R0_BUF_0 (.A(clk_L1_B365), .X(clk_L0_B5841));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R0_INV_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y54__R1_BUF_0 (.A(clk_L1_B367), .X(clk_L0_B5877));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R1_INV_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R2_INV_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R2_INV_1 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y54__R3_BUF_0 (.A(clk_L1_B369), .X(clk_L0_B5913));
  sky130_fd_sc_hd__clkbuf_4 T9Y55__R0_BUF_0 (.A(clk_L1_B371), .X(clk_L0_B5949));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R0_INV_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y55__R1_BUF_0 (.A(clk_L1_B374), .X(clk_L0_B5985));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R1_INV_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R2_INV_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R2_INV_1 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y55__R3_BUF_0 (.A(clk_L1_B376), .X(clk_L0_B6021));
  sky130_fd_sc_hd__clkbuf_4 T9Y56__R0_BUF_0 (.A(clk_L1_B378), .X(clk_L0_B6057));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R0_INV_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y56__R1_BUF_0 (.A(clk_L1_B380), .X(clk_L0_B6093));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R1_INV_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R2_INV_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R2_INV_1 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y56__R3_BUF_0 (.A(clk_L1_B383), .X(clk_L0_B6129));
  sky130_fd_sc_hd__clkbuf_4 T9Y57__R0_BUF_0 (.A(clk_L1_B385), .X(clk_L0_B6165));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R0_INV_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y57__R1_BUF_0 (.A(clk_L1_B387), .X(clk_L0_B6201));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R1_INV_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R2_INV_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R2_INV_1 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y57__R3_BUF_0 (.A(clk_L1_B389), .X(clk_L0_B6237));
  sky130_fd_sc_hd__clkbuf_4 T9Y58__R0_BUF_0 (.A(clk_L1_B392), .X(clk_L0_B6273));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R0_INV_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y58__R1_BUF_0 (.A(clk_L1_B394), .X(clk_L0_B6309));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R1_INV_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R2_INV_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R2_INV_1 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y58__R3_BUF_0 (.A(clk_L1_B396), .X(clk_L0_B6345));
  sky130_fd_sc_hd__clkbuf_4 T9Y59__R0_BUF_0 (.A(clk_L1_B398), .X(clk_L0_B6381));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R0_INV_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y59__R1_BUF_0 (.A(clk_L1_B401), .X(clk_L0_B6417));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R1_INV_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R2_INV_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R2_INV_1 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y59__R3_BUF_0 (.A(clk_L1_B403), .X(clk_L0_B6453));
  sky130_fd_sc_hd__clkbuf_4 T9Y5__R0_BUF_0 (.A(clk_L1_B34), .X(clk_L0_B550));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R0_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y5__R1_BUF_0 (.A(clk_L1_B36), .X(clk_L0_B586));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R1_INV_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R2_INV_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R2_INV_1 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y5__R3_BUF_0 (.A(clk_L1_B38), .X(clk_L0_B622));
  sky130_fd_sc_hd__clkbuf_4 T9Y60__R0_BUF_0 (.A(clk_L1_B405), .X(clk_L0_B6489));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R0_INV_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y60__R1_BUF_0 (.A(clk_L1_B407), .X(clk_L0_B6525));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R1_INV_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R2_INV_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R2_INV_1 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y60__R3_BUF_0 (.A(clk_L1_B410), .X(clk_L0_B6561));
  sky130_fd_sc_hd__clkbuf_4 T9Y61__R0_BUF_0 (.A(clk_L1_B412), .X(clk_L0_B6597));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R0_INV_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y61__R1_BUF_0 (.A(clk_L1_B414), .X(clk_L0_B6633));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R1_INV_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R2_INV_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R2_INV_1 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y61__R3_BUF_0 (.A(clk_L1_B416), .X(clk_L0_B6669));
  sky130_fd_sc_hd__clkbuf_4 T9Y62__R0_BUF_0 (.A(clk_L1_B419), .X(clk_L0_B6705));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R0_INV_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y62__R1_BUF_0 (.A(clk_L1_B421), .X(clk_L0_B6741));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R1_INV_0 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R2_INV_0 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R2_INV_1 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y62__R3_BUF_0 (.A(clk_L1_B423), .X(clk_L0_B6777));
  sky130_fd_sc_hd__clkbuf_4 T9Y63__R0_BUF_0 (.A(clk_L1_B425), .X(clk_L0_B6813));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R0_INV_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y63__R1_BUF_0 (.A(clk_L1_B428), .X(clk_L0_B6849));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R1_INV_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R2_INV_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R2_INV_1 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y63__R3_BUF_0 (.A(clk_L1_B430), .X(clk_L0_B6885));
  sky130_fd_sc_hd__clkbuf_4 T9Y64__R0_BUF_0 (.A(clk_L1_B432), .X(clk_L0_B6921));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R0_INV_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y64__R1_BUF_0 (.A(clk_L1_B434), .X(clk_L0_B6957));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R1_INV_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R2_INV_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R2_INV_1 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y64__R3_BUF_0 (.A(clk_L1_B437), .X(clk_L0_B6993));
  sky130_fd_sc_hd__clkbuf_4 T9Y65__R0_BUF_0 (.A(clk_L1_B439), .X(clk_L0_B7029));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R0_INV_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y65__R1_BUF_0 (.A(clk_L1_B441), .X(clk_L0_B7065));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R1_INV_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R2_INV_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R2_INV_1 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y65__R3_BUF_0 (.A(clk_L1_B443), .X(clk_L0_B7101));
  sky130_fd_sc_hd__clkbuf_4 T9Y66__R0_BUF_0 (.A(clk_L1_B446), .X(clk_L0_B7137));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R0_INV_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y66__R1_BUF_0 (.A(clk_L1_B448), .X(clk_L0_B7173));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R1_INV_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R2_INV_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R2_INV_1 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y66__R3_BUF_0 (.A(clk_L1_B450), .X(clk_L0_B7209));
  sky130_fd_sc_hd__clkbuf_4 T9Y67__R0_BUF_0 (.A(clk_L1_B452), .X(clk_L0_B7245));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R0_INV_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y67__R1_BUF_0 (.A(clk_L1_B455), .X(clk_L0_B7281));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R1_INV_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R2_INV_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R2_INV_1 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y67__R3_BUF_0 (.A(clk_L1_B457), .X(clk_L0_B7317));
  sky130_fd_sc_hd__clkbuf_4 T9Y68__R0_BUF_0 (.A(clk_L1_B459), .X(clk_L0_B7353));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R0_INV_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y68__R1_BUF_0 (.A(clk_L1_B461), .X(clk_L0_B7389));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R1_INV_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R2_INV_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R2_INV_1 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y68__R3_BUF_0 (.A(clk_L1_B464), .X(clk_L0_B7425));
  sky130_fd_sc_hd__clkbuf_4 T9Y69__R0_BUF_0 (.A(clk_L1_B466), .X(clk_L0_B7461));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R0_INV_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y69__R1_BUF_0 (.A(clk_L1_B468), .X(clk_L0_B7497));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R1_INV_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R2_INV_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R2_INV_1 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y69__R3_BUF_0 (.A(clk_L1_B470), .X(clk_L0_B7533));
  sky130_fd_sc_hd__clkbuf_4 T9Y6__R0_BUF_0 (.A(clk_L1_B41), .X(clk_L0_B658));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R0_INV_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y6__R1_BUF_0 (.A(clk_L1_B43), .X(clk_L0_B694));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R1_INV_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R2_INV_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R2_INV_1 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y6__R3_BUF_0 (.A(clk_L1_B45), .X(clk_L0_B730));
  sky130_fd_sc_hd__clkbuf_4 T9Y70__R0_BUF_0 (.A(clk_L1_B473), .X(clk_L0_B7569));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R0_INV_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y70__R1_BUF_0 (.A(clk_L1_B475), .X(clk_L0_B7605));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R1_INV_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R2_INV_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R2_INV_1 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y70__R3_BUF_0 (.A(clk_L1_B477), .X(clk_L0_B7641));
  sky130_fd_sc_hd__clkbuf_4 T9Y71__R0_BUF_0 (.A(clk_L1_B479), .X(clk_L0_B7677));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R0_INV_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y71__R1_BUF_0 (.A(clk_L1_B482), .X(clk_L0_B7713));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R1_INV_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R2_INV_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R2_INV_1 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y71__R3_BUF_0 (.A(clk_L1_B484), .X(clk_L0_B7749));
  sky130_fd_sc_hd__clkbuf_4 T9Y72__R0_BUF_0 (.A(clk_L1_B486), .X(clk_L0_B7785));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R0_INV_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y72__R1_BUF_0 (.A(clk_L1_B488), .X(clk_L0_B7821));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R1_INV_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R2_INV_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R2_INV_1 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y72__R3_BUF_0 (.A(clk_L1_B491), .X(clk_L0_B7857));
  sky130_fd_sc_hd__clkbuf_4 T9Y73__R0_BUF_0 (.A(clk_L1_B493), .X(clk_L0_B7893));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R0_INV_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y73__R1_BUF_0 (.A(clk_L1_B495), .X(clk_L0_B7929));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R1_INV_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R2_INV_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R2_INV_1 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y73__R3_BUF_0 (.A(clk_L1_B497), .X(clk_L0_B7965));
  sky130_fd_sc_hd__clkbuf_4 T9Y74__R0_BUF_0 (.A(clk_L1_B500), .X(clk_L0_B8001));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R0_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y74__R1_BUF_0 (.A(clk_L1_B502), .X(clk_L0_B8037));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R1_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R2_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R2_INV_1 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y74__R3_BUF_0 (.A(clk_L1_B504), .X(clk_L0_B8073));
  sky130_fd_sc_hd__clkbuf_4 T9Y75__R0_BUF_0 (.A(clk_L1_B506), .X(clk_L0_B8109));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R0_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y75__R1_BUF_0 (.A(clk_L1_B509), .X(clk_L0_B8145));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R1_INV_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R2_INV_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R2_INV_1 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y75__R3_BUF_0 (.A(clk_L1_B511), .X(clk_L0_B8181));
  sky130_fd_sc_hd__clkbuf_4 T9Y76__R0_BUF_0 (.A(clk_L1_B513), .X(clk_L0_B8217));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R0_INV_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y76__R1_BUF_0 (.A(clk_L1_B515), .X(clk_L0_B8253));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R1_INV_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R2_INV_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R2_INV_1 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y76__R3_BUF_0 (.A(clk_L1_B518), .X(clk_L0_B8289));
  sky130_fd_sc_hd__clkbuf_4 T9Y77__R0_BUF_0 (.A(clk_L1_B520), .X(clk_L0_B8325));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R0_INV_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y77__R1_BUF_0 (.A(clk_L1_B522), .X(clk_L0_B8361));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R1_INV_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R2_INV_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R2_INV_1 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y77__R3_BUF_0 (.A(clk_L1_B524), .X(clk_L0_B8397));
  sky130_fd_sc_hd__clkbuf_4 T9Y78__R0_BUF_0 (.A(clk_L1_B527), .X(clk_L0_B8433));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R0_INV_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y78__R1_BUF_0 (.A(clk_L1_B529), .X(clk_L0_B8469));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R1_INV_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R2_INV_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R2_INV_1 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y78__R3_BUF_0 (.A(clk_L1_B531), .X(clk_L0_B8505));
  sky130_fd_sc_hd__clkbuf_4 T9Y79__R0_BUF_0 (.A(clk_L1_B533), .X(clk_L0_B8541));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R0_INV_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y79__R1_BUF_0 (.A(clk_L1_B536), .X(clk_L0_B8577));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R1_INV_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R2_INV_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R2_INV_1 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y79__R3_BUF_0 (.A(clk_L1_B538), .X(clk_L0_B8613));
  sky130_fd_sc_hd__clkbuf_4 T9Y7__R0_BUF_0 (.A(clk_L1_B47), .X(clk_L0_B766));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R0_INV_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y7__R1_BUF_0 (.A(clk_L1_B50), .X(clk_L0_B802));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R1_INV_0 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R2_INV_0 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R2_INV_1 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y7__R3_BUF_0 (.A(clk_L1_B52), .X(clk_L0_B838));
  sky130_fd_sc_hd__clkbuf_4 T9Y80__R0_BUF_0 (.A(clk_L1_B540), .X(clk_L0_B8649));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R0_INV_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y80__R1_BUF_0 (.A(clk_L1_B542), .X(clk_L0_B8685));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R1_INV_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R2_INV_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R2_INV_1 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y80__R3_BUF_0 (.A(clk_L1_B545), .X(clk_L0_B8721));
  sky130_fd_sc_hd__clkbuf_4 T9Y81__R0_BUF_0 (.A(clk_L1_B547), .X(clk_L0_B8757));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R0_INV_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y81__R1_BUF_0 (.A(clk_L1_B549), .X(clk_L0_B8793));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R1_INV_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R2_INV_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R2_INV_1 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y81__R3_BUF_0 (.A(clk_L1_B551), .X(clk_L0_B8829));
  sky130_fd_sc_hd__clkbuf_4 T9Y82__R0_BUF_0 (.A(clk_L1_B554), .X(clk_L0_B8865));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R0_INV_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y82__R1_BUF_0 (.A(clk_L1_B556), .X(clk_L0_B8901));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R1_INV_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R2_INV_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R2_INV_1 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y82__R3_BUF_0 (.A(clk_L1_B558), .X(clk_L0_B8937));
  sky130_fd_sc_hd__clkbuf_4 T9Y83__R0_BUF_0 (.A(clk_L1_B560), .X(clk_L0_B8973));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R0_INV_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y83__R1_BUF_0 (.A(clk_L1_B563), .X(clk_L0_B9009));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R1_INV_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R2_INV_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R2_INV_1 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y83__R3_BUF_0 (.A(clk_L1_B565), .X(clk_L0_B9045));
  sky130_fd_sc_hd__clkbuf_4 T9Y84__R0_BUF_0 (.A(clk_L1_B567), .X(clk_L0_B9081));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R0_INV_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y84__R1_BUF_0 (.A(clk_L1_B569), .X(clk_L0_B9117));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R1_INV_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R2_INV_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R2_INV_1 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y84__R3_BUF_0 (.A(clk_L1_B572), .X(clk_L0_B9153));
  sky130_fd_sc_hd__clkbuf_4 T9Y85__R0_BUF_0 (.A(clk_L1_B574), .X(clk_L0_B9189));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R0_INV_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y85__R1_BUF_0 (.A(clk_L1_B576), .X(clk_L0_B9225));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R1_INV_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R2_INV_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R2_INV_1 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y85__R3_BUF_0 (.A(clk_L1_B578), .X(clk_L0_B9261));
  sky130_fd_sc_hd__clkbuf_4 T9Y86__R0_BUF_0 (.A(clk_L1_B581), .X(clk_L0_B9297));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R0_INV_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y86__R1_BUF_0 (.A(clk_L1_B583), .X(clk_L0_B9333));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R1_INV_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R2_INV_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R2_INV_1 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y86__R3_BUF_0 (.A(clk_L1_B585), .X(clk_L0_B9369));
  sky130_fd_sc_hd__clkbuf_4 T9Y87__R0_BUF_0 (.A(clk_L1_B587), .X(clk_L0_B9405));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R0_INV_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y87__R1_BUF_0 (.A(clk_L1_B590), .X(clk_L0_B9441));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R1_INV_0 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R2_INV_0 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R2_INV_1 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y87__R3_BUF_0 (.A(clk_L1_B592), .X(clk_L0_B9477));
  sky130_fd_sc_hd__clkbuf_4 T9Y88__R0_BUF_0 (.A(clk_L1_B594), .X(clk_L0_B9513));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R0_INV_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y88__R1_BUF_0 (.A(clk_L1_B596), .X(clk_L0_B9549));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R1_INV_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R2_INV_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R2_INV_1 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y88__R3_BUF_0 (.A(clk_L1_B599), .X(clk_L0_B9585));
  sky130_fd_sc_hd__clkbuf_4 T9Y89__R0_BUF_0 (.A(clk_L1_B601), .X(clk_L0_B9621));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R0_INV_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y89__R1_BUF_0 (.A(clk_L1_B603), .X(clk_L0_B9657));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R1_INV_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R2_INV_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R2_INV_1 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y89__R3_BUF_0 (.A(clk_L1_B605), .X(clk_L0_B9693));
  sky130_fd_sc_hd__clkbuf_4 T9Y8__R0_BUF_0 (.A(clk_L1_B54), .X(clk_L0_B874));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R0_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y8__R1_BUF_0 (.A(clk_L1_B56), .X(clk_L0_B910));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R1_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R2_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R2_INV_1 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y8__R3_BUF_0 (.A(clk_L1_B59), .X(clk_L0_B946));
  sky130_fd_sc_hd__clkbuf_4 T9Y9__R0_BUF_0 (.A(clk_L1_B61), .X(clk_L0_B982));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R0_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y9__R1_BUF_0 (.A(clk_L1_B63), .X(clk_L0_B1018));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R1_INV_0 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R2_INV_0 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R2_INV_1 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y9__R3_BUF_0 (.A(clk_L1_B65), .X(clk_L0_B1054));

endmodule
