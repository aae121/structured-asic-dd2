// 6502 Final Netlist with CTS and ECO
// Design cells: 28819
// CTS/ECO cells: 0
// Total: 28819

module 6502_final (clk, rst_n, in_0, in_1, in_2, in_3, in_4, in_5, in_6, in_7, in_8, in_9, in_10, in_11, in_12, in_13, in_14, in_15, in_16, in_17, in_18, in_19, in_20, in_21, in_22, in_23, in_24, in_25, in_26, in_27, in_28, in_29, in_30, in_31, in_32, in_33, in_34, in_35, in_36, in_37, in_38, in_39, oeb_0, oeb_1, oeb_2, oeb_3, oeb_4, oeb_5, oeb_6, oeb_7, oeb_8, oeb_9, oeb_10, oeb_11, oeb_12, oeb_13, oeb_14, oeb_15, oeb_16, oeb_17, oeb_18, oeb_19, oeb_20, oeb_21, oeb_22, oeb_23, oeb_24, oeb_25, oeb_26, oeb_27, oeb_28, oeb_29, oeb_30, oeb_31, oeb_32, oeb_33, oeb_34, oeb_35, oeb_36, oeb_37, oeb_38, oeb_39, out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21, out_22, out_23, out_24, out_25, out_26, out_27, out_28, out_29, out_30, out_31, out_32, out_33, out_34, out_35, out_36, out_37, out_38, out_39);

  input clk;
  input rst_n;
  input in_0;
  input in_1;
  input in_2;
  input in_3;
  input in_4;
  input in_5;
  input in_6;
  input in_7;
  input in_8;
  input in_9;
  input in_10;
  input in_11;
  input in_12;
  input in_13;
  input in_14;
  input in_15;
  input in_16;
  input in_17;
  input in_18;
  input in_19;
  input in_20;
  input in_21;
  input in_22;
  input in_23;
  input in_24;
  input in_25;
  input in_26;
  input in_27;
  input in_28;
  input in_29;
  input in_30;
  input in_31;
  input in_32;
  input in_33;
  input in_34;
  input in_35;
  input in_36;
  input in_37;
  input in_38;
  input in_39;
  output oeb_0;
  output oeb_1;
  output oeb_2;
  output oeb_3;
  output oeb_4;
  output oeb_5;
  output oeb_6;
  output oeb_7;
  output oeb_8;
  output oeb_9;
  output oeb_10;
  output oeb_11;
  output oeb_12;
  output oeb_13;
  output oeb_14;
  output oeb_15;
  output oeb_16;
  output oeb_17;
  output oeb_18;
  output oeb_19;
  output oeb_20;
  output oeb_21;
  output oeb_22;
  output oeb_23;
  output oeb_24;
  output oeb_25;
  output oeb_26;
  output oeb_27;
  output oeb_28;
  output oeb_29;
  output oeb_30;
  output oeb_31;
  output oeb_32;
  output oeb_33;
  output oeb_34;
  output oeb_35;
  output oeb_36;
  output oeb_37;
  output oeb_38;
  output oeb_39;
  output out_0;
  output out_1;
  output out_2;
  output out_3;
  output out_4;
  output out_5;
  output out_6;
  output out_7;
  output out_8;
  output out_9;
  output out_10;
  output out_11;
  output out_12;
  output out_13;
  output out_14;
  output out_15;
  output out_16;
  output out_17;
  output out_18;
  output out_19;
  output out_20;
  output out_21;
  output out_22;
  output out_23;
  output out_24;
  output out_25;
  output out_26;
  output out_27;
  output out_28;
  output out_29;
  output out_30;
  output out_31;
  output out_32;
  output out_33;
  output out_34;
  output out_35;
  output out_36;
  output out_37;
  output out_38;
  output out_39;

  // Internal nets
  wire 100;
  wire 1000;
  wire 1001;
  wire 1002;
  wire 1003;
  wire 1004;
  wire 1005;
  wire 1006;
  wire 1007;
  wire 1008;
  wire 1009;
  wire 101;
  wire 1010;
  wire 1011;
  wire 1012;
  wire 1013;
  wire 1014;
  wire 1015;
  wire 1016;
  wire 1017;
  wire 1018;
  wire 1019;
  wire 102;
  wire 1020;
  wire 1021;
  wire 1022;
  wire 1023;
  wire 1024;
  wire 1025;
  wire 1026;
  wire 1027;
  wire 1028;
  wire 1029;
  wire 103;
  wire 1030;
  wire 1031;
  wire 1032;
  wire 1033;
  wire 1034;
  wire 1035;
  wire 1036;
  wire 1037;
  wire 1038;
  wire 1039;
  wire 104;
  wire 1040;
  wire 1041;
  wire 1042;
  wire 1043;
  wire 1044;
  wire 1045;
  wire 1046;
  wire 1047;
  wire 1048;
  wire 1049;
  wire 105;
  wire 1050;
  wire 1051;
  wire 1052;
  wire 1053;
  wire 1054;
  wire 1055;
  wire 1056;
  wire 1057;
  wire 1058;
  wire 1059;
  wire 106;
  wire 1060;
  wire 1061;
  wire 1062;
  wire 1063;
  wire 1064;
  wire 1065;
  wire 1066;
  wire 1067;
  wire 1068;
  wire 1069;
  wire 107;
  wire 1070;
  wire 1071;
  wire 1072;
  wire 1073;
  wire 1074;
  wire 1075;
  wire 1076;
  wire 1077;
  wire 1078;
  wire 1079;
  wire 108;
  wire 1080;
  wire 1081;
  wire 1082;
  wire 1083;
  wire 1084;
  wire 1085;
  wire 1086;
  wire 1087;
  wire 1088;
  wire 1089;
  wire 109;
  wire 1090;
  wire 1091;
  wire 1092;
  wire 1093;
  wire 1094;
  wire 1095;
  wire 1096;
  wire 1097;
  wire 1098;
  wire 1099;
  wire 110;
  wire 1100;
  wire 1101;
  wire 1102;
  wire 1103;
  wire 1104;
  wire 1105;
  wire 1106;
  wire 1107;
  wire 1108;
  wire 1109;
  wire 111;
  wire 1110;
  wire 1111;
  wire 1112;
  wire 1113;
  wire 1114;
  wire 1115;
  wire 1116;
  wire 1117;
  wire 1118;
  wire 1119;
  wire 112;
  wire 1120;
  wire 1121;
  wire 1122;
  wire 1123;
  wire 1124;
  wire 1125;
  wire 1126;
  wire 1127;
  wire 1128;
  wire 1129;
  wire 113;
  wire 1130;
  wire 1131;
  wire 1132;
  wire 1133;
  wire 1134;
  wire 1135;
  wire 1136;
  wire 1137;
  wire 1138;
  wire 1139;
  wire 114;
  wire 1140;
  wire 1141;
  wire 1142;
  wire 1143;
  wire 1144;
  wire 1145;
  wire 1146;
  wire 1147;
  wire 1148;
  wire 1149;
  wire 115;
  wire 1150;
  wire 1151;
  wire 1152;
  wire 1153;
  wire 1154;
  wire 1155;
  wire 1156;
  wire 1157;
  wire 1158;
  wire 1159;
  wire 116;
  wire 1160;
  wire 1161;
  wire 1162;
  wire 1163;
  wire 1164;
  wire 1165;
  wire 1166;
  wire 1167;
  wire 1168;
  wire 1169;
  wire 117;
  wire 1170;
  wire 1171;
  wire 1172;
  wire 1173;
  wire 1174;
  wire 1175;
  wire 1176;
  wire 1177;
  wire 1178;
  wire 1179;
  wire 118;
  wire 1180;
  wire 1181;
  wire 1182;
  wire 1183;
  wire 1184;
  wire 1185;
  wire 1186;
  wire 1187;
  wire 1188;
  wire 1189;
  wire 119;
  wire 1190;
  wire 1191;
  wire 1192;
  wire 1193;
  wire 1194;
  wire 1195;
  wire 1196;
  wire 1197;
  wire 1198;
  wire 1199;
  wire 120;
  wire 1200;
  wire 1201;
  wire 1202;
  wire 1203;
  wire 1204;
  wire 1205;
  wire 1206;
  wire 1207;
  wire 1208;
  wire 1209;
  wire 121;
  wire 1210;
  wire 1211;
  wire 1212;
  wire 1213;
  wire 1214;
  wire 1215;
  wire 1216;
  wire 1217;
  wire 1218;
  wire 1219;
  wire 122;
  wire 1220;
  wire 1221;
  wire 1222;
  wire 1223;
  wire 1224;
  wire 1225;
  wire 1226;
  wire 1227;
  wire 1228;
  wire 1229;
  wire 123;
  wire 1230;
  wire 1231;
  wire 1232;
  wire 1233;
  wire 1234;
  wire 1235;
  wire 1236;
  wire 1237;
  wire 1238;
  wire 1239;
  wire 124;
  wire 1240;
  wire 1241;
  wire 1242;
  wire 1243;
  wire 1244;
  wire 1245;
  wire 1246;
  wire 1247;
  wire 1248;
  wire 1249;
  wire 125;
  wire 1250;
  wire 1251;
  wire 1252;
  wire 1253;
  wire 1254;
  wire 1255;
  wire 1256;
  wire 1257;
  wire 1258;
  wire 1259;
  wire 126;
  wire 1260;
  wire 1261;
  wire 1262;
  wire 1263;
  wire 1264;
  wire 1265;
  wire 1266;
  wire 1267;
  wire 1268;
  wire 1269;
  wire 127;
  wire 1270;
  wire 1271;
  wire 1272;
  wire 1273;
  wire 1274;
  wire 1275;
  wire 1276;
  wire 1277;
  wire 1278;
  wire 1279;
  wire 128;
  wire 1280;
  wire 1281;
  wire 1282;
  wire 1283;
  wire 1284;
  wire 1285;
  wire 1286;
  wire 1287;
  wire 1288;
  wire 1289;
  wire 129;
  wire 1290;
  wire 1291;
  wire 1292;
  wire 1293;
  wire 1294;
  wire 1295;
  wire 1296;
  wire 1297;
  wire 1298;
  wire 1299;
  wire 130;
  wire 1300;
  wire 1301;
  wire 1302;
  wire 1303;
  wire 1304;
  wire 1305;
  wire 1306;
  wire 1307;
  wire 1308;
  wire 1309;
  wire 131;
  wire 1310;
  wire 1311;
  wire 1312;
  wire 1313;
  wire 1314;
  wire 1315;
  wire 1316;
  wire 1317;
  wire 1318;
  wire 1319;
  wire 132;
  wire 1320;
  wire 1321;
  wire 1322;
  wire 1323;
  wire 1324;
  wire 1325;
  wire 1326;
  wire 1327;
  wire 1328;
  wire 1329;
  wire 133;
  wire 1330;
  wire 1331;
  wire 1332;
  wire 1333;
  wire 1334;
  wire 1335;
  wire 1336;
  wire 1337;
  wire 1338;
  wire 1339;
  wire 134;
  wire 1340;
  wire 1341;
  wire 1342;
  wire 1343;
  wire 1344;
  wire 1345;
  wire 1346;
  wire 1347;
  wire 1348;
  wire 1349;
  wire 135;
  wire 1350;
  wire 1351;
  wire 1352;
  wire 1353;
  wire 1354;
  wire 1355;
  wire 1356;
  wire 1357;
  wire 1358;
  wire 1359;
  wire 136;
  wire 1360;
  wire 1361;
  wire 1362;
  wire 1363;
  wire 1364;
  wire 1365;
  wire 1366;
  wire 1367;
  wire 1368;
  wire 1369;
  wire 137;
  wire 1370;
  wire 1371;
  wire 1372;
  wire 1373;
  wire 1374;
  wire 1375;
  wire 1376;
  wire 1377;
  wire 1378;
  wire 1379;
  wire 138;
  wire 1380;
  wire 1381;
  wire 1382;
  wire 1383;
  wire 1384;
  wire 1385;
  wire 1386;
  wire 1387;
  wire 1388;
  wire 1389;
  wire 139;
  wire 1390;
  wire 1391;
  wire 1392;
  wire 1393;
  wire 1394;
  wire 1395;
  wire 1396;
  wire 1397;
  wire 1398;
  wire 1399;
  wire 140;
  wire 1400;
  wire 1401;
  wire 1402;
  wire 1403;
  wire 1404;
  wire 1405;
  wire 1406;
  wire 1407;
  wire 1408;
  wire 1409;
  wire 141;
  wire 1410;
  wire 1411;
  wire 1412;
  wire 1413;
  wire 1414;
  wire 1415;
  wire 1416;
  wire 1417;
  wire 1418;
  wire 1419;
  wire 142;
  wire 1420;
  wire 1421;
  wire 1422;
  wire 1423;
  wire 1424;
  wire 1425;
  wire 1426;
  wire 1427;
  wire 1428;
  wire 1429;
  wire 143;
  wire 1430;
  wire 1431;
  wire 1432;
  wire 1433;
  wire 1434;
  wire 1435;
  wire 1436;
  wire 1437;
  wire 1438;
  wire 1439;
  wire 144;
  wire 1440;
  wire 1441;
  wire 1442;
  wire 1443;
  wire 1444;
  wire 1445;
  wire 1446;
  wire 1447;
  wire 1448;
  wire 1449;
  wire 145;
  wire 1450;
  wire 1451;
  wire 1452;
  wire 1453;
  wire 1454;
  wire 1455;
  wire 1456;
  wire 1457;
  wire 1458;
  wire 1459;
  wire 146;
  wire 1460;
  wire 1461;
  wire 1462;
  wire 1463;
  wire 1464;
  wire 1465;
  wire 1466;
  wire 1467;
  wire 1468;
  wire 1469;
  wire 147;
  wire 1470;
  wire 1471;
  wire 1472;
  wire 1473;
  wire 1474;
  wire 1475;
  wire 1476;
  wire 1477;
  wire 1478;
  wire 1479;
  wire 148;
  wire 1480;
  wire 1481;
  wire 1482;
  wire 1483;
  wire 1484;
  wire 1485;
  wire 1486;
  wire 1487;
  wire 1488;
  wire 1489;
  wire 149;
  wire 1490;
  wire 1491;
  wire 1492;
  wire 1493;
  wire 1494;
  wire 1495;
  wire 1496;
  wire 1497;
  wire 1498;
  wire 1499;
  wire 150;
  wire 1500;
  wire 1501;
  wire 1502;
  wire 1503;
  wire 1504;
  wire 1505;
  wire 1506;
  wire 1507;
  wire 1508;
  wire 1509;
  wire 151;
  wire 1510;
  wire 1511;
  wire 1512;
  wire 1513;
  wire 1514;
  wire 1515;
  wire 1516;
  wire 1517;
  wire 1518;
  wire 1519;
  wire 152;
  wire 1520;
  wire 1521;
  wire 1522;
  wire 1523;
  wire 1524;
  wire 1525;
  wire 1526;
  wire 1527;
  wire 1528;
  wire 1529;
  wire 153;
  wire 1530;
  wire 1531;
  wire 1532;
  wire 1533;
  wire 1534;
  wire 1535;
  wire 1536;
  wire 1537;
  wire 1538;
  wire 1539;
  wire 154;
  wire 1540;
  wire 1541;
  wire 1542;
  wire 1543;
  wire 1544;
  wire 1545;
  wire 1546;
  wire 1547;
  wire 1548;
  wire 1549;
  wire 155;
  wire 1550;
  wire 1551;
  wire 1552;
  wire 1553;
  wire 1554;
  wire 1555;
  wire 1556;
  wire 1557;
  wire 1558;
  wire 1559;
  wire 156;
  wire 1560;
  wire 1561;
  wire 1562;
  wire 1563;
  wire 1564;
  wire 1565;
  wire 1566;
  wire 1567;
  wire 1568;
  wire 1569;
  wire 157;
  wire 1570;
  wire 1571;
  wire 1572;
  wire 1573;
  wire 1574;
  wire 1575;
  wire 1576;
  wire 1577;
  wire 1578;
  wire 1579;
  wire 158;
  wire 1580;
  wire 1581;
  wire 1582;
  wire 1583;
  wire 1584;
  wire 1585;
  wire 1586;
  wire 1587;
  wire 1588;
  wire 1589;
  wire 159;
  wire 1590;
  wire 1591;
  wire 1592;
  wire 1593;
  wire 1594;
  wire 1595;
  wire 1596;
  wire 1597;
  wire 1598;
  wire 1599;
  wire 160;
  wire 1600;
  wire 1601;
  wire 1602;
  wire 1603;
  wire 1604;
  wire 1605;
  wire 1606;
  wire 1607;
  wire 1608;
  wire 1609;
  wire 161;
  wire 1610;
  wire 1611;
  wire 1612;
  wire 1613;
  wire 1614;
  wire 1615;
  wire 1616;
  wire 1617;
  wire 1618;
  wire 1619;
  wire 162;
  wire 1620;
  wire 1621;
  wire 1622;
  wire 1623;
  wire 1624;
  wire 1625;
  wire 1626;
  wire 1627;
  wire 1628;
  wire 1629;
  wire 163;
  wire 1630;
  wire 1631;
  wire 1632;
  wire 1633;
  wire 1634;
  wire 1635;
  wire 1636;
  wire 1637;
  wire 1638;
  wire 1639;
  wire 164;
  wire 1640;
  wire 1641;
  wire 1642;
  wire 1643;
  wire 1644;
  wire 1645;
  wire 1646;
  wire 1647;
  wire 1648;
  wire 1649;
  wire 165;
  wire 1650;
  wire 1651;
  wire 1652;
  wire 1653;
  wire 1654;
  wire 1655;
  wire 1656;
  wire 1657;
  wire 1658;
  wire 1659;
  wire 166;
  wire 1660;
  wire 1661;
  wire 1662;
  wire 1663;
  wire 1664;
  wire 1665;
  wire 1666;
  wire 1667;
  wire 1668;
  wire 1669;
  wire 167;
  wire 1670;
  wire 1671;
  wire 1672;
  wire 1673;
  wire 1674;
  wire 1675;
  wire 1676;
  wire 1677;
  wire 1678;
  wire 1679;
  wire 168;
  wire 1680;
  wire 1681;
  wire 1682;
  wire 1683;
  wire 1684;
  wire 1685;
  wire 1686;
  wire 1687;
  wire 1688;
  wire 1689;
  wire 169;
  wire 1690;
  wire 1691;
  wire 1692;
  wire 1693;
  wire 1694;
  wire 1695;
  wire 1696;
  wire 1697;
  wire 1698;
  wire 1699;
  wire 170;
  wire 1700;
  wire 1701;
  wire 1702;
  wire 1703;
  wire 1704;
  wire 1705;
  wire 1706;
  wire 1707;
  wire 1708;
  wire 1709;
  wire 171;
  wire 1710;
  wire 1711;
  wire 1712;
  wire 1713;
  wire 1714;
  wire 1715;
  wire 1716;
  wire 1717;
  wire 1718;
  wire 1719;
  wire 172;
  wire 1720;
  wire 1721;
  wire 1722;
  wire 1723;
  wire 1724;
  wire 1725;
  wire 1726;
  wire 1727;
  wire 1728;
  wire 1729;
  wire 173;
  wire 1730;
  wire 1731;
  wire 1732;
  wire 1733;
  wire 1734;
  wire 1735;
  wire 1736;
  wire 1737;
  wire 1738;
  wire 1739;
  wire 174;
  wire 1740;
  wire 1741;
  wire 1742;
  wire 1743;
  wire 1744;
  wire 1745;
  wire 1746;
  wire 1747;
  wire 1748;
  wire 1749;
  wire 175;
  wire 1750;
  wire 1751;
  wire 1752;
  wire 1753;
  wire 1754;
  wire 1755;
  wire 1756;
  wire 1757;
  wire 1758;
  wire 1759;
  wire 176;
  wire 1760;
  wire 1761;
  wire 1762;
  wire 1763;
  wire 1764;
  wire 1765;
  wire 1766;
  wire 1767;
  wire 1768;
  wire 1769;
  wire 177;
  wire 1770;
  wire 1771;
  wire 1772;
  wire 1773;
  wire 1774;
  wire 1775;
  wire 1776;
  wire 1777;
  wire 1778;
  wire 1779;
  wire 178;
  wire 1780;
  wire 1781;
  wire 1782;
  wire 1783;
  wire 1784;
  wire 1785;
  wire 1786;
  wire 1787;
  wire 1788;
  wire 1789;
  wire 179;
  wire 1790;
  wire 1791;
  wire 1792;
  wire 1793;
  wire 1794;
  wire 1795;
  wire 1796;
  wire 1797;
  wire 1798;
  wire 1799;
  wire 180;
  wire 1800;
  wire 1801;
  wire 1802;
  wire 1803;
  wire 1804;
  wire 1805;
  wire 1806;
  wire 1807;
  wire 1808;
  wire 1809;
  wire 181;
  wire 1810;
  wire 1811;
  wire 1812;
  wire 1813;
  wire 1814;
  wire 1815;
  wire 1816;
  wire 1817;
  wire 1818;
  wire 1819;
  wire 182;
  wire 1820;
  wire 1821;
  wire 1822;
  wire 1823;
  wire 1824;
  wire 1825;
  wire 1826;
  wire 1827;
  wire 1828;
  wire 1829;
  wire 183;
  wire 1830;
  wire 1831;
  wire 1832;
  wire 1833;
  wire 1834;
  wire 1835;
  wire 1836;
  wire 1837;
  wire 1838;
  wire 1839;
  wire 184;
  wire 1840;
  wire 1841;
  wire 1842;
  wire 1843;
  wire 1844;
  wire 1845;
  wire 1846;
  wire 1847;
  wire 1848;
  wire 1849;
  wire 185;
  wire 1850;
  wire 1851;
  wire 1852;
  wire 1853;
  wire 1854;
  wire 1855;
  wire 1856;
  wire 1857;
  wire 1858;
  wire 1859;
  wire 186;
  wire 1860;
  wire 1861;
  wire 1862;
  wire 1863;
  wire 1864;
  wire 1865;
  wire 1866;
  wire 1867;
  wire 1868;
  wire 1869;
  wire 187;
  wire 1870;
  wire 1871;
  wire 1872;
  wire 1873;
  wire 1874;
  wire 1875;
  wire 1876;
  wire 1877;
  wire 1878;
  wire 1879;
  wire 188;
  wire 1880;
  wire 1881;
  wire 1882;
  wire 1883;
  wire 1884;
  wire 1885;
  wire 1886;
  wire 1887;
  wire 1888;
  wire 1889;
  wire 189;
  wire 1890;
  wire 1891;
  wire 1892;
  wire 1893;
  wire 1894;
  wire 1895;
  wire 1896;
  wire 1897;
  wire 1898;
  wire 1899;
  wire 190;
  wire 1900;
  wire 1901;
  wire 1902;
  wire 1903;
  wire 1904;
  wire 1905;
  wire 1906;
  wire 1907;
  wire 1908;
  wire 1909;
  wire 191;
  wire 1910;
  wire 1911;
  wire 1912;
  wire 1913;
  wire 1914;
  wire 1915;
  wire 1916;
  wire 1917;
  wire 1918;
  wire 1919;
  wire 192;
  wire 1920;
  wire 1921;
  wire 1922;
  wire 1923;
  wire 1924;
  wire 1925;
  wire 1926;
  wire 1927;
  wire 1928;
  wire 1929;
  wire 193;
  wire 1930;
  wire 1931;
  wire 1932;
  wire 1933;
  wire 1934;
  wire 1935;
  wire 1936;
  wire 1937;
  wire 1938;
  wire 1939;
  wire 194;
  wire 1940;
  wire 1941;
  wire 1942;
  wire 1943;
  wire 1944;
  wire 1945;
  wire 1946;
  wire 1947;
  wire 1948;
  wire 1949;
  wire 195;
  wire 1950;
  wire 1951;
  wire 1952;
  wire 1953;
  wire 1954;
  wire 1955;
  wire 1956;
  wire 1957;
  wire 1958;
  wire 1959;
  wire 196;
  wire 1960;
  wire 1961;
  wire 1962;
  wire 1963;
  wire 1964;
  wire 1965;
  wire 1966;
  wire 1967;
  wire 1968;
  wire 1969;
  wire 197;
  wire 1970;
  wire 1971;
  wire 1972;
  wire 1973;
  wire 1974;
  wire 1975;
  wire 1976;
  wire 1977;
  wire 1978;
  wire 1979;
  wire 198;
  wire 1980;
  wire 1981;
  wire 1982;
  wire 1983;
  wire 1984;
  wire 1985;
  wire 1986;
  wire 1987;
  wire 1988;
  wire 1989;
  wire 199;
  wire 1990;
  wire 1991;
  wire 1992;
  wire 1993;
  wire 1994;
  wire 1995;
  wire 1996;
  wire 1997;
  wire 1998;
  wire 1999;
  wire 2;
  wire 20;
  wire 200;
  wire 2000;
  wire 2001;
  wire 2002;
  wire 2003;
  wire 2004;
  wire 2005;
  wire 2006;
  wire 2007;
  wire 2008;
  wire 2009;
  wire 201;
  wire 2010;
  wire 2011;
  wire 2012;
  wire 2013;
  wire 2014;
  wire 2015;
  wire 2016;
  wire 2017;
  wire 2018;
  wire 2019;
  wire 202;
  wire 2020;
  wire 2021;
  wire 2022;
  wire 2023;
  wire 2024;
  wire 2025;
  wire 2026;
  wire 2027;
  wire 2028;
  wire 2029;
  wire 203;
  wire 2030;
  wire 2031;
  wire 2032;
  wire 2033;
  wire 2034;
  wire 2035;
  wire 2036;
  wire 2037;
  wire 2038;
  wire 2039;
  wire 204;
  wire 2040;
  wire 2041;
  wire 2042;
  wire 2043;
  wire 2044;
  wire 2045;
  wire 2046;
  wire 2047;
  wire 2048;
  wire 2049;
  wire 205;
  wire 2050;
  wire 2051;
  wire 2052;
  wire 2053;
  wire 2054;
  wire 2055;
  wire 2056;
  wire 2057;
  wire 2058;
  wire 2059;
  wire 206;
  wire 2060;
  wire 2061;
  wire 2062;
  wire 2063;
  wire 2064;
  wire 2065;
  wire 2066;
  wire 2067;
  wire 2068;
  wire 2069;
  wire 207;
  wire 2070;
  wire 2071;
  wire 2072;
  wire 2073;
  wire 2074;
  wire 2075;
  wire 2076;
  wire 2077;
  wire 2078;
  wire 2079;
  wire 208;
  wire 2080;
  wire 2081;
  wire 2082;
  wire 2083;
  wire 2084;
  wire 2085;
  wire 2086;
  wire 2087;
  wire 2088;
  wire 2089;
  wire 209;
  wire 2090;
  wire 2091;
  wire 2092;
  wire 2093;
  wire 2094;
  wire 2095;
  wire 2096;
  wire 2097;
  wire 2098;
  wire 2099;
  wire 21;
  wire 210;
  wire 2100;
  wire 2101;
  wire 2102;
  wire 2103;
  wire 2104;
  wire 2105;
  wire 2106;
  wire 2107;
  wire 2108;
  wire 2109;
  wire 211;
  wire 2110;
  wire 2111;
  wire 2112;
  wire 2113;
  wire 2114;
  wire 2115;
  wire 2116;
  wire 2117;
  wire 2118;
  wire 2119;
  wire 212;
  wire 2120;
  wire 2121;
  wire 2122;
  wire 2123;
  wire 2124;
  wire 2125;
  wire 2126;
  wire 2127;
  wire 2128;
  wire 2129;
  wire 213;
  wire 2130;
  wire 2131;
  wire 2132;
  wire 2133;
  wire 2134;
  wire 2135;
  wire 2136;
  wire 2137;
  wire 2138;
  wire 2139;
  wire 214;
  wire 2140;
  wire 2141;
  wire 2142;
  wire 2143;
  wire 2144;
  wire 2145;
  wire 2146;
  wire 2147;
  wire 2148;
  wire 2149;
  wire 215;
  wire 2150;
  wire 2151;
  wire 2152;
  wire 2153;
  wire 2154;
  wire 2155;
  wire 2156;
  wire 2157;
  wire 2158;
  wire 2159;
  wire 216;
  wire 2160;
  wire 2161;
  wire 2162;
  wire 2163;
  wire 2164;
  wire 2165;
  wire 2166;
  wire 2167;
  wire 2168;
  wire 2169;
  wire 217;
  wire 2170;
  wire 2171;
  wire 2172;
  wire 2173;
  wire 2174;
  wire 2175;
  wire 2176;
  wire 2177;
  wire 2178;
  wire 2179;
  wire 218;
  wire 2180;
  wire 2181;
  wire 2182;
  wire 2183;
  wire 2184;
  wire 2185;
  wire 2186;
  wire 2187;
  wire 2188;
  wire 2189;
  wire 219;
  wire 2190;
  wire 2191;
  wire 2192;
  wire 2193;
  wire 2194;
  wire 2195;
  wire 2196;
  wire 2197;
  wire 2198;
  wire 2199;
  wire 22;
  wire 220;
  wire 2200;
  wire 2201;
  wire 2202;
  wire 2203;
  wire 2204;
  wire 2205;
  wire 2206;
  wire 2207;
  wire 2208;
  wire 2209;
  wire 221;
  wire 2210;
  wire 2211;
  wire 2212;
  wire 2213;
  wire 2214;
  wire 2215;
  wire 2216;
  wire 2217;
  wire 2218;
  wire 2219;
  wire 222;
  wire 2220;
  wire 2221;
  wire 2222;
  wire 2223;
  wire 2224;
  wire 2225;
  wire 2226;
  wire 2227;
  wire 2228;
  wire 2229;
  wire 223;
  wire 2230;
  wire 2231;
  wire 2232;
  wire 2233;
  wire 2234;
  wire 2235;
  wire 2236;
  wire 2237;
  wire 2238;
  wire 2239;
  wire 224;
  wire 2240;
  wire 2241;
  wire 2242;
  wire 2243;
  wire 2244;
  wire 2245;
  wire 2246;
  wire 2247;
  wire 2248;
  wire 2249;
  wire 225;
  wire 2250;
  wire 2251;
  wire 2252;
  wire 2253;
  wire 2254;
  wire 2255;
  wire 2256;
  wire 2257;
  wire 2258;
  wire 2259;
  wire 226;
  wire 2260;
  wire 2261;
  wire 2262;
  wire 2263;
  wire 2264;
  wire 2265;
  wire 2266;
  wire 2267;
  wire 2268;
  wire 2269;
  wire 227;
  wire 2270;
  wire 2271;
  wire 2272;
  wire 2273;
  wire 2274;
  wire 2275;
  wire 2276;
  wire 2277;
  wire 2278;
  wire 2279;
  wire 228;
  wire 2280;
  wire 2281;
  wire 2282;
  wire 2283;
  wire 2284;
  wire 2285;
  wire 2286;
  wire 2287;
  wire 2288;
  wire 2289;
  wire 229;
  wire 2290;
  wire 2291;
  wire 2292;
  wire 2293;
  wire 2294;
  wire 2295;
  wire 2296;
  wire 2297;
  wire 2298;
  wire 2299;
  wire 23;
  wire 230;
  wire 2300;
  wire 2301;
  wire 2302;
  wire 2303;
  wire 2304;
  wire 2305;
  wire 2306;
  wire 2307;
  wire 2308;
  wire 2309;
  wire 231;
  wire 2310;
  wire 2311;
  wire 2312;
  wire 2313;
  wire 2314;
  wire 2315;
  wire 2316;
  wire 2317;
  wire 2318;
  wire 2319;
  wire 232;
  wire 2320;
  wire 2321;
  wire 2322;
  wire 2323;
  wire 2324;
  wire 2325;
  wire 2326;
  wire 2327;
  wire 2328;
  wire 2329;
  wire 233;
  wire 2330;
  wire 2331;
  wire 2332;
  wire 2333;
  wire 2334;
  wire 2335;
  wire 2336;
  wire 2337;
  wire 2338;
  wire 2339;
  wire 234;
  wire 2340;
  wire 2341;
  wire 2342;
  wire 2343;
  wire 2344;
  wire 2345;
  wire 2346;
  wire 2347;
  wire 2348;
  wire 2349;
  wire 235;
  wire 2350;
  wire 2351;
  wire 2352;
  wire 2353;
  wire 2354;
  wire 2355;
  wire 2356;
  wire 2357;
  wire 2358;
  wire 2359;
  wire 236;
  wire 2360;
  wire 2361;
  wire 2362;
  wire 2363;
  wire 2364;
  wire 2365;
  wire 2366;
  wire 2367;
  wire 2368;
  wire 2369;
  wire 237;
  wire 2370;
  wire 2371;
  wire 2372;
  wire 2373;
  wire 2374;
  wire 2375;
  wire 2376;
  wire 2377;
  wire 2378;
  wire 2379;
  wire 238;
  wire 2380;
  wire 2381;
  wire 2382;
  wire 2383;
  wire 2384;
  wire 2385;
  wire 2386;
  wire 2387;
  wire 2388;
  wire 2389;
  wire 239;
  wire 2390;
  wire 2391;
  wire 2392;
  wire 2393;
  wire 2394;
  wire 2395;
  wire 2396;
  wire 2397;
  wire 2398;
  wire 2399;
  wire 24;
  wire 240;
  wire 2400;
  wire 2401;
  wire 2402;
  wire 2403;
  wire 2404;
  wire 2405;
  wire 2406;
  wire 2407;
  wire 2408;
  wire 2409;
  wire 241;
  wire 2410;
  wire 2411;
  wire 2412;
  wire 2413;
  wire 2414;
  wire 2415;
  wire 2416;
  wire 2417;
  wire 2418;
  wire 2419;
  wire 242;
  wire 2420;
  wire 2421;
  wire 2422;
  wire 2423;
  wire 2424;
  wire 2425;
  wire 2426;
  wire 2427;
  wire 2428;
  wire 2429;
  wire 243;
  wire 2430;
  wire 2431;
  wire 2432;
  wire 2433;
  wire 2434;
  wire 2435;
  wire 2436;
  wire 2437;
  wire 2438;
  wire 2439;
  wire 244;
  wire 2440;
  wire 2441;
  wire 2442;
  wire 2443;
  wire 2444;
  wire 2445;
  wire 2446;
  wire 2447;
  wire 2448;
  wire 2449;
  wire 245;
  wire 2450;
  wire 2451;
  wire 2452;
  wire 2453;
  wire 2454;
  wire 2455;
  wire 2456;
  wire 2457;
  wire 2458;
  wire 2459;
  wire 246;
  wire 2460;
  wire 2461;
  wire 2462;
  wire 2463;
  wire 2464;
  wire 2465;
  wire 2466;
  wire 2467;
  wire 2468;
  wire 2469;
  wire 247;
  wire 2470;
  wire 2471;
  wire 2472;
  wire 2473;
  wire 2474;
  wire 2475;
  wire 2476;
  wire 2477;
  wire 2478;
  wire 2479;
  wire 248;
  wire 2480;
  wire 2481;
  wire 2482;
  wire 2483;
  wire 2484;
  wire 2485;
  wire 2486;
  wire 2487;
  wire 2488;
  wire 2489;
  wire 249;
  wire 2490;
  wire 2491;
  wire 2492;
  wire 2493;
  wire 2494;
  wire 2495;
  wire 2496;
  wire 2497;
  wire 2498;
  wire 2499;
  wire 25;
  wire 250;
  wire 2500;
  wire 2501;
  wire 2502;
  wire 2503;
  wire 2504;
  wire 2505;
  wire 2506;
  wire 2507;
  wire 2508;
  wire 2509;
  wire 251;
  wire 2510;
  wire 2511;
  wire 2512;
  wire 2513;
  wire 2514;
  wire 2515;
  wire 2516;
  wire 2517;
  wire 2518;
  wire 2519;
  wire 252;
  wire 2520;
  wire 2521;
  wire 2522;
  wire 2523;
  wire 2524;
  wire 2525;
  wire 2526;
  wire 2527;
  wire 2528;
  wire 2529;
  wire 253;
  wire 2530;
  wire 2531;
  wire 2532;
  wire 2533;
  wire 2534;
  wire 2535;
  wire 2536;
  wire 2537;
  wire 2538;
  wire 2539;
  wire 254;
  wire 2540;
  wire 2541;
  wire 2542;
  wire 2543;
  wire 2544;
  wire 2545;
  wire 2546;
  wire 2547;
  wire 2548;
  wire 2549;
  wire 255;
  wire 2550;
  wire 2551;
  wire 2552;
  wire 2553;
  wire 2554;
  wire 2555;
  wire 2556;
  wire 2557;
  wire 2558;
  wire 2559;
  wire 256;
  wire 2560;
  wire 2561;
  wire 2562;
  wire 2563;
  wire 2564;
  wire 2565;
  wire 2566;
  wire 2567;
  wire 2568;
  wire 2569;
  wire 257;
  wire 2570;
  wire 2571;
  wire 2572;
  wire 2573;
  wire 2574;
  wire 2575;
  wire 2576;
  wire 2577;
  wire 2578;
  wire 2579;
  wire 258;
  wire 2580;
  wire 2581;
  wire 2582;
  wire 2583;
  wire 2584;
  wire 2585;
  wire 2586;
  wire 2587;
  wire 2588;
  wire 2589;
  wire 259;
  wire 2590;
  wire 2591;
  wire 2592;
  wire 2593;
  wire 2594;
  wire 2595;
  wire 2596;
  wire 2597;
  wire 2598;
  wire 2599;
  wire 26;
  wire 260;
  wire 2600;
  wire 2601;
  wire 2602;
  wire 2603;
  wire 2604;
  wire 2605;
  wire 2606;
  wire 2607;
  wire 2608;
  wire 2609;
  wire 261;
  wire 2610;
  wire 2611;
  wire 2612;
  wire 2613;
  wire 2614;
  wire 2615;
  wire 2616;
  wire 2617;
  wire 2618;
  wire 2619;
  wire 262;
  wire 2620;
  wire 2621;
  wire 2622;
  wire 2623;
  wire 2624;
  wire 2625;
  wire 2626;
  wire 2627;
  wire 2628;
  wire 2629;
  wire 263;
  wire 2630;
  wire 2631;
  wire 2632;
  wire 2633;
  wire 2634;
  wire 2635;
  wire 2636;
  wire 2637;
  wire 2638;
  wire 2639;
  wire 264;
  wire 2640;
  wire 2641;
  wire 2642;
  wire 2643;
  wire 2644;
  wire 2645;
  wire 2646;
  wire 2647;
  wire 2648;
  wire 2649;
  wire 265;
  wire 2650;
  wire 2651;
  wire 2652;
  wire 2653;
  wire 2654;
  wire 2655;
  wire 2656;
  wire 2657;
  wire 2658;
  wire 2659;
  wire 266;
  wire 2660;
  wire 2661;
  wire 2662;
  wire 2663;
  wire 2664;
  wire 2665;
  wire 2666;
  wire 2667;
  wire 2668;
  wire 2669;
  wire 267;
  wire 2670;
  wire 2671;
  wire 2672;
  wire 2673;
  wire 2674;
  wire 2675;
  wire 2676;
  wire 2677;
  wire 2678;
  wire 2679;
  wire 268;
  wire 2680;
  wire 2681;
  wire 2682;
  wire 2683;
  wire 2684;
  wire 2685;
  wire 2686;
  wire 2687;
  wire 2688;
  wire 2689;
  wire 269;
  wire 2690;
  wire 2691;
  wire 2692;
  wire 2693;
  wire 2694;
  wire 2695;
  wire 2696;
  wire 2697;
  wire 2698;
  wire 2699;
  wire 27;
  wire 270;
  wire 2700;
  wire 2701;
  wire 2702;
  wire 2703;
  wire 2704;
  wire 2705;
  wire 2706;
  wire 2707;
  wire 2708;
  wire 2709;
  wire 271;
  wire 2710;
  wire 2711;
  wire 2712;
  wire 2713;
  wire 2714;
  wire 2715;
  wire 2716;
  wire 2717;
  wire 2718;
  wire 2719;
  wire 272;
  wire 2720;
  wire 2721;
  wire 2722;
  wire 2723;
  wire 2724;
  wire 2725;
  wire 2726;
  wire 2727;
  wire 2728;
  wire 2729;
  wire 273;
  wire 2730;
  wire 2731;
  wire 2732;
  wire 2733;
  wire 2734;
  wire 2735;
  wire 2736;
  wire 2737;
  wire 2738;
  wire 2739;
  wire 274;
  wire 2740;
  wire 2741;
  wire 2742;
  wire 2743;
  wire 2744;
  wire 2745;
  wire 2746;
  wire 2747;
  wire 2748;
  wire 2749;
  wire 275;
  wire 2750;
  wire 2751;
  wire 2752;
  wire 2753;
  wire 2754;
  wire 2755;
  wire 2756;
  wire 2757;
  wire 2758;
  wire 2759;
  wire 276;
  wire 2760;
  wire 2761;
  wire 2762;
  wire 2763;
  wire 2764;
  wire 2765;
  wire 2766;
  wire 2767;
  wire 2768;
  wire 2769;
  wire 277;
  wire 2770;
  wire 2771;
  wire 2772;
  wire 2773;
  wire 2774;
  wire 2775;
  wire 2776;
  wire 2777;
  wire 2778;
  wire 2779;
  wire 278;
  wire 2780;
  wire 2781;
  wire 2782;
  wire 2783;
  wire 2784;
  wire 2785;
  wire 2786;
  wire 2787;
  wire 2788;
  wire 2789;
  wire 279;
  wire 2790;
  wire 2791;
  wire 2792;
  wire 2793;
  wire 2794;
  wire 2795;
  wire 2796;
  wire 2797;
  wire 2798;
  wire 2799;
  wire 280;
  wire 2800;
  wire 2801;
  wire 2802;
  wire 2803;
  wire 2804;
  wire 2805;
  wire 2806;
  wire 2807;
  wire 2808;
  wire 2809;
  wire 281;
  wire 2810;
  wire 2811;
  wire 2812;
  wire 2813;
  wire 2814;
  wire 2815;
  wire 2816;
  wire 2817;
  wire 2818;
  wire 2819;
  wire 282;
  wire 2820;
  wire 2821;
  wire 2822;
  wire 2823;
  wire 2824;
  wire 2825;
  wire 2826;
  wire 2827;
  wire 2828;
  wire 2829;
  wire 283;
  wire 2830;
  wire 2831;
  wire 2832;
  wire 2833;
  wire 2834;
  wire 2835;
  wire 2836;
  wire 2837;
  wire 2838;
  wire 2839;
  wire 284;
  wire 2840;
  wire 2841;
  wire 2842;
  wire 2843;
  wire 2844;
  wire 2845;
  wire 2846;
  wire 2847;
  wire 2848;
  wire 2849;
  wire 285;
  wire 2850;
  wire 2851;
  wire 2852;
  wire 2853;
  wire 2854;
  wire 2855;
  wire 2856;
  wire 2857;
  wire 2858;
  wire 2859;
  wire 286;
  wire 2860;
  wire 2861;
  wire 2862;
  wire 2863;
  wire 2864;
  wire 2865;
  wire 2866;
  wire 2867;
  wire 2868;
  wire 2869;
  wire 287;
  wire 2870;
  wire 2871;
  wire 2872;
  wire 2873;
  wire 2874;
  wire 2875;
  wire 2876;
  wire 2877;
  wire 2878;
  wire 2879;
  wire 288;
  wire 2880;
  wire 2881;
  wire 2882;
  wire 2883;
  wire 2884;
  wire 2885;
  wire 2886;
  wire 2887;
  wire 2888;
  wire 2889;
  wire 289;
  wire 2890;
  wire 2891;
  wire 2892;
  wire 2893;
  wire 2894;
  wire 2895;
  wire 2896;
  wire 2897;
  wire 2898;
  wire 2899;
  wire 290;
  wire 2900;
  wire 2901;
  wire 2902;
  wire 2903;
  wire 2904;
  wire 2905;
  wire 2906;
  wire 2907;
  wire 2908;
  wire 2909;
  wire 291;
  wire 2910;
  wire 2911;
  wire 2912;
  wire 2913;
  wire 2914;
  wire 2915;
  wire 2916;
  wire 2917;
  wire 2918;
  wire 2919;
  wire 292;
  wire 2920;
  wire 2921;
  wire 2922;
  wire 2923;
  wire 2924;
  wire 2925;
  wire 2926;
  wire 2927;
  wire 2928;
  wire 2929;
  wire 293;
  wire 2930;
  wire 2931;
  wire 2932;
  wire 2933;
  wire 2934;
  wire 2935;
  wire 2936;
  wire 2937;
  wire 2938;
  wire 2939;
  wire 294;
  wire 2940;
  wire 2941;
  wire 2942;
  wire 2943;
  wire 2944;
  wire 2945;
  wire 2946;
  wire 2947;
  wire 2948;
  wire 2949;
  wire 295;
  wire 2950;
  wire 2951;
  wire 2952;
  wire 2953;
  wire 2954;
  wire 2955;
  wire 2956;
  wire 2957;
  wire 2958;
  wire 2959;
  wire 296;
  wire 2960;
  wire 2961;
  wire 2962;
  wire 2963;
  wire 2964;
  wire 2965;
  wire 2966;
  wire 2967;
  wire 2968;
  wire 2969;
  wire 297;
  wire 2970;
  wire 2971;
  wire 2972;
  wire 2973;
  wire 2974;
  wire 2975;
  wire 2976;
  wire 2977;
  wire 2978;
  wire 2979;
  wire 298;
  wire 2980;
  wire 2981;
  wire 2982;
  wire 2983;
  wire 2984;
  wire 2985;
  wire 2986;
  wire 2987;
  wire 2988;
  wire 2989;
  wire 299;
  wire 2990;
  wire 2991;
  wire 2992;
  wire 2993;
  wire 2994;
  wire 2995;
  wire 2996;
  wire 2997;
  wire 2998;
  wire 2999;
  wire 3;
  wire 300;
  wire 3000;
  wire 3001;
  wire 3002;
  wire 3003;
  wire 3004;
  wire 3005;
  wire 3006;
  wire 3007;
  wire 3008;
  wire 3009;
  wire 301;
  wire 3010;
  wire 3011;
  wire 3012;
  wire 3013;
  wire 3014;
  wire 3015;
  wire 3016;
  wire 3017;
  wire 3018;
  wire 3019;
  wire 302;
  wire 3020;
  wire 3021;
  wire 3022;
  wire 3023;
  wire 3024;
  wire 3025;
  wire 3026;
  wire 3027;
  wire 3028;
  wire 3029;
  wire 303;
  wire 3030;
  wire 3031;
  wire 3032;
  wire 3033;
  wire 3034;
  wire 3035;
  wire 3036;
  wire 3037;
  wire 3038;
  wire 3039;
  wire 304;
  wire 3040;
  wire 3041;
  wire 3042;
  wire 3043;
  wire 3044;
  wire 3045;
  wire 3046;
  wire 3047;
  wire 3048;
  wire 3049;
  wire 305;
  wire 3050;
  wire 3051;
  wire 3052;
  wire 3053;
  wire 3054;
  wire 3055;
  wire 3056;
  wire 3057;
  wire 3058;
  wire 3059;
  wire 306;
  wire 3060;
  wire 3061;
  wire 3062;
  wire 3063;
  wire 3064;
  wire 3065;
  wire 3066;
  wire 3067;
  wire 3068;
  wire 3069;
  wire 307;
  wire 3070;
  wire 3071;
  wire 3072;
  wire 3073;
  wire 3074;
  wire 3075;
  wire 3076;
  wire 3077;
  wire 3078;
  wire 3079;
  wire 308;
  wire 3080;
  wire 3081;
  wire 3082;
  wire 3083;
  wire 3084;
  wire 3085;
  wire 3086;
  wire 3087;
  wire 309;
  wire 310;
  wire 311;
  wire 312;
  wire 313;
  wire 314;
  wire 315;
  wire 316;
  wire 317;
  wire 318;
  wire 319;
  wire 320;
  wire 321;
  wire 322;
  wire 323;
  wire 324;
  wire 325;
  wire 326;
  wire 327;
  wire 328;
  wire 329;
  wire 330;
  wire 331;
  wire 332;
  wire 333;
  wire 334;
  wire 335;
  wire 336;
  wire 337;
  wire 338;
  wire 339;
  wire 340;
  wire 341;
  wire 342;
  wire 343;
  wire 344;
  wire 345;
  wire 346;
  wire 347;
  wire 348;
  wire 349;
  wire 350;
  wire 351;
  wire 352;
  wire 353;
  wire 354;
  wire 355;
  wire 356;
  wire 357;
  wire 358;
  wire 359;
  wire 360;
  wire 361;
  wire 362;
  wire 363;
  wire 364;
  wire 365;
  wire 366;
  wire 367;
  wire 368;
  wire 369;
  wire 37;
  wire 370;
  wire 371;
  wire 372;
  wire 373;
  wire 374;
  wire 375;
  wire 376;
  wire 377;
  wire 378;
  wire 379;
  wire 38;
  wire 380;
  wire 381;
  wire 382;
  wire 383;
  wire 384;
  wire 385;
  wire 386;
  wire 387;
  wire 388;
  wire 389;
  wire 39;
  wire 390;
  wire 391;
  wire 392;
  wire 393;
  wire 394;
  wire 395;
  wire 396;
  wire 397;
  wire 398;
  wire 399;
  wire 400;
  wire 401;
  wire 402;
  wire 403;
  wire 404;
  wire 405;
  wire 406;
  wire 407;
  wire 408;
  wire 409;
  wire 410;
  wire 411;
  wire 412;
  wire 413;
  wire 414;
  wire 415;
  wire 416;
  wire 417;
  wire 418;
  wire 419;
  wire 420;
  wire 421;
  wire 422;
  wire 423;
  wire 424;
  wire 425;
  wire 426;
  wire 427;
  wire 428;
  wire 429;
  wire 430;
  wire 431;
  wire 432;
  wire 433;
  wire 434;
  wire 435;
  wire 436;
  wire 437;
  wire 438;
  wire 439;
  wire 44;
  wire 440;
  wire 441;
  wire 442;
  wire 443;
  wire 444;
  wire 445;
  wire 446;
  wire 447;
  wire 448;
  wire 449;
  wire 45;
  wire 450;
  wire 451;
  wire 452;
  wire 453;
  wire 454;
  wire 455;
  wire 456;
  wire 457;
  wire 458;
  wire 459;
  wire 46;
  wire 460;
  wire 461;
  wire 462;
  wire 463;
  wire 464;
  wire 465;
  wire 466;
  wire 467;
  wire 468;
  wire 469;
  wire 47;
  wire 470;
  wire 471;
  wire 472;
  wire 473;
  wire 474;
  wire 475;
  wire 476;
  wire 477;
  wire 478;
  wire 479;
  wire 48;
  wire 480;
  wire 481;
  wire 482;
  wire 483;
  wire 484;
  wire 485;
  wire 486;
  wire 487;
  wire 488;
  wire 489;
  wire 49;
  wire 490;
  wire 491;
  wire 492;
  wire 493;
  wire 494;
  wire 495;
  wire 496;
  wire 497;
  wire 498;
  wire 499;
  wire 50;
  wire 500;
  wire 501;
  wire 502;
  wire 503;
  wire 504;
  wire 505;
  wire 506;
  wire 507;
  wire 508;
  wire 509;
  wire 51;
  wire 510;
  wire 511;
  wire 512;
  wire 513;
  wire 514;
  wire 515;
  wire 516;
  wire 517;
  wire 518;
  wire 519;
  wire 52;
  wire 520;
  wire 521;
  wire 522;
  wire 523;
  wire 524;
  wire 525;
  wire 526;
  wire 527;
  wire 528;
  wire 529;
  wire 53;
  wire 530;
  wire 531;
  wire 532;
  wire 533;
  wire 534;
  wire 535;
  wire 536;
  wire 537;
  wire 538;
  wire 539;
  wire 54;
  wire 540;
  wire 541;
  wire 542;
  wire 543;
  wire 544;
  wire 545;
  wire 546;
  wire 547;
  wire 548;
  wire 549;
  wire 55;
  wire 550;
  wire 551;
  wire 552;
  wire 553;
  wire 554;
  wire 555;
  wire 556;
  wire 557;
  wire 558;
  wire 559;
  wire 56;
  wire 560;
  wire 561;
  wire 562;
  wire 563;
  wire 564;
  wire 565;
  wire 566;
  wire 567;
  wire 568;
  wire 569;
  wire 57;
  wire 570;
  wire 571;
  wire 572;
  wire 573;
  wire 574;
  wire 575;
  wire 576;
  wire 577;
  wire 578;
  wire 579;
  wire 58;
  wire 580;
  wire 581;
  wire 582;
  wire 583;
  wire 584;
  wire 585;
  wire 586;
  wire 587;
  wire 588;
  wire 589;
  wire 59;
  wire 590;
  wire 591;
  wire 592;
  wire 593;
  wire 594;
  wire 595;
  wire 596;
  wire 597;
  wire 598;
  wire 599;
  wire 60;
  wire 600;
  wire 601;
  wire 602;
  wire 603;
  wire 604;
  wire 605;
  wire 606;
  wire 607;
  wire 608;
  wire 609;
  wire 61;
  wire 610;
  wire 611;
  wire 612;
  wire 613;
  wire 614;
  wire 615;
  wire 616;
  wire 617;
  wire 618;
  wire 619;
  wire 62;
  wire 620;
  wire 621;
  wire 622;
  wire 623;
  wire 624;
  wire 625;
  wire 626;
  wire 627;
  wire 628;
  wire 629;
  wire 63;
  wire 630;
  wire 631;
  wire 632;
  wire 633;
  wire 634;
  wire 635;
  wire 636;
  wire 637;
  wire 638;
  wire 639;
  wire 64;
  wire 640;
  wire 641;
  wire 642;
  wire 643;
  wire 644;
  wire 645;
  wire 646;
  wire 647;
  wire 648;
  wire 649;
  wire 65;
  wire 650;
  wire 651;
  wire 652;
  wire 653;
  wire 654;
  wire 655;
  wire 656;
  wire 657;
  wire 658;
  wire 659;
  wire 66;
  wire 660;
  wire 661;
  wire 662;
  wire 663;
  wire 664;
  wire 665;
  wire 666;
  wire 667;
  wire 668;
  wire 669;
  wire 67;
  wire 670;
  wire 671;
  wire 672;
  wire 673;
  wire 674;
  wire 675;
  wire 676;
  wire 677;
  wire 678;
  wire 679;
  wire 68;
  wire 680;
  wire 681;
  wire 682;
  wire 683;
  wire 684;
  wire 685;
  wire 686;
  wire 687;
  wire 688;
  wire 689;
  wire 69;
  wire 690;
  wire 691;
  wire 692;
  wire 693;
  wire 694;
  wire 695;
  wire 696;
  wire 697;
  wire 698;
  wire 699;
  wire 70;
  wire 700;
  wire 701;
  wire 702;
  wire 703;
  wire 704;
  wire 705;
  wire 706;
  wire 707;
  wire 708;
  wire 709;
  wire 71;
  wire 710;
  wire 711;
  wire 712;
  wire 713;
  wire 714;
  wire 715;
  wire 716;
  wire 717;
  wire 718;
  wire 719;
  wire 72;
  wire 720;
  wire 721;
  wire 722;
  wire 723;
  wire 724;
  wire 725;
  wire 726;
  wire 727;
  wire 728;
  wire 729;
  wire 73;
  wire 730;
  wire 731;
  wire 732;
  wire 733;
  wire 734;
  wire 735;
  wire 736;
  wire 737;
  wire 738;
  wire 739;
  wire 74;
  wire 740;
  wire 741;
  wire 742;
  wire 743;
  wire 744;
  wire 745;
  wire 746;
  wire 747;
  wire 748;
  wire 749;
  wire 75;
  wire 750;
  wire 751;
  wire 752;
  wire 753;
  wire 754;
  wire 755;
  wire 756;
  wire 757;
  wire 758;
  wire 759;
  wire 76;
  wire 760;
  wire 761;
  wire 762;
  wire 763;
  wire 764;
  wire 765;
  wire 766;
  wire 767;
  wire 768;
  wire 769;
  wire 77;
  wire 770;
  wire 771;
  wire 772;
  wire 773;
  wire 774;
  wire 775;
  wire 776;
  wire 777;
  wire 778;
  wire 779;
  wire 78;
  wire 780;
  wire 781;
  wire 782;
  wire 783;
  wire 784;
  wire 785;
  wire 786;
  wire 787;
  wire 788;
  wire 789;
  wire 79;
  wire 790;
  wire 791;
  wire 792;
  wire 793;
  wire 794;
  wire 795;
  wire 796;
  wire 797;
  wire 798;
  wire 799;
  wire 80;
  wire 800;
  wire 801;
  wire 802;
  wire 803;
  wire 804;
  wire 805;
  wire 806;
  wire 807;
  wire 808;
  wire 809;
  wire 81;
  wire 810;
  wire 811;
  wire 812;
  wire 813;
  wire 814;
  wire 815;
  wire 816;
  wire 817;
  wire 818;
  wire 819;
  wire 82;
  wire 820;
  wire 821;
  wire 822;
  wire 823;
  wire 824;
  wire 825;
  wire 826;
  wire 827;
  wire 828;
  wire 829;
  wire 83;
  wire 830;
  wire 831;
  wire 832;
  wire 833;
  wire 834;
  wire 835;
  wire 836;
  wire 837;
  wire 838;
  wire 839;
  wire 84;
  wire 840;
  wire 841;
  wire 842;
  wire 843;
  wire 844;
  wire 845;
  wire 846;
  wire 847;
  wire 848;
  wire 849;
  wire 85;
  wire 850;
  wire 851;
  wire 852;
  wire 853;
  wire 854;
  wire 855;
  wire 856;
  wire 857;
  wire 858;
  wire 859;
  wire 86;
  wire 860;
  wire 861;
  wire 862;
  wire 863;
  wire 864;
  wire 865;
  wire 866;
  wire 867;
  wire 868;
  wire 869;
  wire 87;
  wire 870;
  wire 871;
  wire 872;
  wire 873;
  wire 874;
  wire 875;
  wire 876;
  wire 877;
  wire 878;
  wire 879;
  wire 88;
  wire 880;
  wire 881;
  wire 882;
  wire 883;
  wire 884;
  wire 885;
  wire 886;
  wire 887;
  wire 888;
  wire 889;
  wire 89;
  wire 890;
  wire 891;
  wire 892;
  wire 893;
  wire 894;
  wire 895;
  wire 896;
  wire 897;
  wire 898;
  wire 899;
  wire 90;
  wire 900;
  wire 901;
  wire 902;
  wire 903;
  wire 904;
  wire 905;
  wire 906;
  wire 907;
  wire 908;
  wire 909;
  wire 91;
  wire 910;
  wire 911;
  wire 912;
  wire 913;
  wire 914;
  wire 915;
  wire 916;
  wire 917;
  wire 918;
  wire 919;
  wire 92;
  wire 920;
  wire 921;
  wire 922;
  wire 923;
  wire 924;
  wire 925;
  wire 926;
  wire 927;
  wire 928;
  wire 929;
  wire 93;
  wire 930;
  wire 931;
  wire 932;
  wire 933;
  wire 934;
  wire 935;
  wire 936;
  wire 937;
  wire 938;
  wire 939;
  wire 94;
  wire 940;
  wire 941;
  wire 942;
  wire 943;
  wire 944;
  wire 945;
  wire 946;
  wire 947;
  wire 948;
  wire 949;
  wire 95;
  wire 950;
  wire 951;
  wire 952;
  wire 953;
  wire 954;
  wire 955;
  wire 956;
  wire 957;
  wire 958;
  wire 959;
  wire 96;
  wire 960;
  wire 961;
  wire 962;
  wire 963;
  wire 964;
  wire 965;
  wire 966;
  wire 967;
  wire 968;
  wire 969;
  wire 97;
  wire 970;
  wire 971;
  wire 972;
  wire 973;
  wire 974;
  wire 975;
  wire 976;
  wire 977;
  wire 978;
  wire 979;
  wire 98;
  wire 980;
  wire 981;
  wire 982;
  wire 983;
  wire 984;
  wire 985;
  wire 986;
  wire 987;
  wire 988;
  wire 989;
  wire 99;
  wire 990;
  wire 991;
  wire 992;
  wire 993;
  wire 994;
  wire 995;
  wire 996;
  wire 997;
  wire 998;
  wire 999;
  wire tie_lo_T0Y0__R2_CONB_0;
  wire tie_lo_T0Y10__R2_CONB_0;
  wire tie_lo_T0Y11__R2_CONB_0;
  wire tie_lo_T0Y12__R2_CONB_0;
  wire tie_lo_T0Y13__R2_CONB_0;
  wire tie_lo_T0Y14__R2_CONB_0;
  wire tie_lo_T0Y15__R2_CONB_0;
  wire tie_lo_T0Y16__R2_CONB_0;
  wire tie_lo_T0Y17__R2_CONB_0;
  wire tie_lo_T0Y18__R2_CONB_0;
  wire tie_lo_T0Y19__R2_CONB_0;
  wire tie_lo_T0Y1__R2_CONB_0;
  wire tie_lo_T0Y20__R2_CONB_0;
  wire tie_lo_T0Y21__R2_CONB_0;
  wire tie_lo_T0Y22__R2_CONB_0;
  wire tie_lo_T0Y23__R2_CONB_0;
  wire tie_lo_T0Y24__R2_CONB_0;
  wire tie_lo_T0Y25__R2_CONB_0;
  wire tie_lo_T0Y26__R2_CONB_0;
  wire tie_lo_T0Y27__R2_CONB_0;
  wire tie_lo_T0Y28__R2_CONB_0;
  wire tie_lo_T0Y29__R2_CONB_0;
  wire tie_lo_T0Y2__R2_CONB_0;
  wire tie_lo_T0Y30__R2_CONB_0;
  wire tie_lo_T0Y31__R2_CONB_0;
  wire tie_lo_T0Y32__R2_CONB_0;
  wire tie_lo_T0Y33__R2_CONB_0;
  wire tie_lo_T0Y34__R2_CONB_0;
  wire tie_lo_T0Y35__R2_CONB_0;
  wire tie_lo_T0Y36__R2_CONB_0;
  wire tie_lo_T0Y37__R2_CONB_0;
  wire tie_lo_T0Y38__R2_CONB_0;
  wire tie_lo_T0Y39__R2_CONB_0;
  wire tie_lo_T0Y3__R2_CONB_0;
  wire tie_lo_T0Y40__R2_CONB_0;
  wire tie_lo_T0Y41__R2_CONB_0;
  wire tie_lo_T0Y42__R2_CONB_0;
  wire tie_lo_T0Y43__R2_CONB_0;
  wire tie_lo_T0Y44__R2_CONB_0;
  wire tie_lo_T0Y45__R2_CONB_0;
  wire tie_lo_T0Y46__R2_CONB_0;
  wire tie_lo_T0Y47__R2_CONB_0;
  wire tie_lo_T0Y48__R2_CONB_0;
  wire tie_lo_T0Y49__R2_CONB_0;
  wire tie_lo_T0Y4__R2_CONB_0;
  wire tie_lo_T0Y50__R2_CONB_0;
  wire tie_lo_T0Y51__R2_CONB_0;
  wire tie_lo_T0Y52__R2_CONB_0;
  wire tie_lo_T0Y53__R2_CONB_0;
  wire tie_lo_T0Y54__R2_CONB_0;
  wire tie_lo_T0Y55__R2_CONB_0;
  wire tie_lo_T0Y56__R2_CONB_0;
  wire tie_lo_T0Y57__R2_CONB_0;
  wire tie_lo_T0Y58__R2_CONB_0;
  wire tie_lo_T0Y59__R2_CONB_0;
  wire tie_lo_T0Y5__R2_CONB_0;
  wire tie_lo_T0Y60__R2_CONB_0;
  wire tie_lo_T0Y61__R2_CONB_0;
  wire tie_lo_T0Y62__R2_CONB_0;
  wire tie_lo_T0Y63__R2_CONB_0;
  wire tie_lo_T0Y64__R2_CONB_0;
  wire tie_lo_T0Y65__R2_CONB_0;
  wire tie_lo_T0Y66__R2_CONB_0;
  wire tie_lo_T0Y67__R2_CONB_0;
  wire tie_lo_T0Y68__R2_CONB_0;
  wire tie_lo_T0Y69__R2_CONB_0;
  wire tie_lo_T0Y6__R2_CONB_0;
  wire tie_lo_T0Y70__R2_CONB_0;
  wire tie_lo_T0Y71__R2_CONB_0;
  wire tie_lo_T0Y72__R2_CONB_0;
  wire tie_lo_T0Y73__R2_CONB_0;
  wire tie_lo_T0Y74__R2_CONB_0;
  wire tie_lo_T0Y75__R2_CONB_0;
  wire tie_lo_T0Y76__R2_CONB_0;
  wire tie_lo_T0Y77__R2_CONB_0;
  wire tie_lo_T0Y78__R2_CONB_0;
  wire tie_lo_T0Y79__R2_CONB_0;
  wire tie_lo_T0Y7__R2_CONB_0;
  wire tie_lo_T0Y80__R2_CONB_0;
  wire tie_lo_T0Y81__R2_CONB_0;
  wire tie_lo_T0Y82__R2_CONB_0;
  wire tie_lo_T0Y83__R2_CONB_0;
  wire tie_lo_T0Y84__R2_CONB_0;
  wire tie_lo_T0Y85__R2_CONB_0;
  wire tie_lo_T0Y86__R2_CONB_0;
  wire tie_lo_T0Y87__R2_CONB_0;
  wire tie_lo_T0Y88__R2_CONB_0;
  wire tie_lo_T0Y89__R2_CONB_0;
  wire tie_lo_T0Y8__R2_CONB_0;
  wire tie_lo_T0Y9__R2_CONB_0;
  wire tie_lo_T10Y0__R2_CONB_0;
  wire tie_lo_T10Y10__R2_CONB_0;
  wire tie_lo_T10Y11__R2_CONB_0;
  wire tie_lo_T10Y12__R2_CONB_0;
  wire tie_lo_T10Y13__R2_CONB_0;
  wire tie_lo_T10Y14__R2_CONB_0;
  wire tie_lo_T10Y15__R2_CONB_0;
  wire tie_lo_T10Y16__R2_CONB_0;
  wire tie_lo_T10Y17__R2_CONB_0;
  wire tie_lo_T10Y18__R2_CONB_0;
  wire tie_lo_T10Y19__R2_CONB_0;
  wire tie_lo_T10Y1__R2_CONB_0;
  wire tie_lo_T10Y20__R2_CONB_0;
  wire tie_lo_T10Y21__R2_CONB_0;
  wire tie_lo_T10Y22__R2_CONB_0;
  wire tie_lo_T10Y23__R2_CONB_0;
  wire tie_lo_T10Y24__R2_CONB_0;
  wire tie_lo_T10Y25__R2_CONB_0;
  wire tie_lo_T10Y26__R2_CONB_0;
  wire tie_lo_T10Y27__R2_CONB_0;
  wire tie_lo_T10Y28__R2_CONB_0;
  wire tie_lo_T10Y29__R2_CONB_0;
  wire tie_lo_T10Y2__R2_CONB_0;
  wire tie_lo_T10Y30__R2_CONB_0;
  wire tie_lo_T10Y31__R2_CONB_0;
  wire tie_lo_T10Y32__R2_CONB_0;
  wire tie_lo_T10Y33__R2_CONB_0;
  wire tie_lo_T10Y34__R2_CONB_0;
  wire tie_lo_T10Y35__R2_CONB_0;
  wire tie_lo_T10Y36__R2_CONB_0;
  wire tie_lo_T10Y37__R2_CONB_0;
  wire tie_lo_T10Y38__R2_CONB_0;
  wire tie_lo_T10Y39__R2_CONB_0;
  wire tie_lo_T10Y3__R2_CONB_0;
  wire tie_lo_T10Y40__R2_CONB_0;
  wire tie_lo_T10Y41__R2_CONB_0;
  wire tie_lo_T10Y42__R2_CONB_0;
  wire tie_lo_T10Y43__R2_CONB_0;
  wire tie_lo_T10Y44__R2_CONB_0;
  wire tie_lo_T10Y45__R2_CONB_0;
  wire tie_lo_T10Y46__R2_CONB_0;
  wire tie_lo_T10Y47__R2_CONB_0;
  wire tie_lo_T10Y48__R2_CONB_0;
  wire tie_lo_T10Y49__R2_CONB_0;
  wire tie_lo_T10Y4__R2_CONB_0;
  wire tie_lo_T10Y50__R2_CONB_0;
  wire tie_lo_T10Y51__R2_CONB_0;
  wire tie_lo_T10Y52__R2_CONB_0;
  wire tie_lo_T10Y53__R2_CONB_0;
  wire tie_lo_T10Y54__R2_CONB_0;
  wire tie_lo_T10Y55__R2_CONB_0;
  wire tie_lo_T10Y56__R2_CONB_0;
  wire tie_lo_T10Y57__R2_CONB_0;
  wire tie_lo_T10Y58__R2_CONB_0;
  wire tie_lo_T10Y59__R2_CONB_0;
  wire tie_lo_T10Y5__R2_CONB_0;
  wire tie_lo_T10Y60__R2_CONB_0;
  wire tie_lo_T10Y61__R2_CONB_0;
  wire tie_lo_T10Y62__R2_CONB_0;
  wire tie_lo_T10Y63__R2_CONB_0;
  wire tie_lo_T10Y64__R2_CONB_0;
  wire tie_lo_T10Y65__R2_CONB_0;
  wire tie_lo_T10Y66__R2_CONB_0;
  wire tie_lo_T10Y67__R2_CONB_0;
  wire tie_lo_T10Y68__R2_CONB_0;
  wire tie_lo_T10Y69__R2_CONB_0;
  wire tie_lo_T10Y6__R2_CONB_0;
  wire tie_lo_T10Y70__R2_CONB_0;
  wire tie_lo_T10Y71__R2_CONB_0;
  wire tie_lo_T10Y72__R2_CONB_0;
  wire tie_lo_T10Y73__R2_CONB_0;
  wire tie_lo_T10Y74__R2_CONB_0;
  wire tie_lo_T10Y75__R2_CONB_0;
  wire tie_lo_T10Y76__R2_CONB_0;
  wire tie_lo_T10Y77__R2_CONB_0;
  wire tie_lo_T10Y78__R2_CONB_0;
  wire tie_lo_T10Y79__R2_CONB_0;
  wire tie_lo_T10Y7__R2_CONB_0;
  wire tie_lo_T10Y80__R2_CONB_0;
  wire tie_lo_T10Y81__R2_CONB_0;
  wire tie_lo_T10Y82__R2_CONB_0;
  wire tie_lo_T10Y83__R2_CONB_0;
  wire tie_lo_T10Y84__R2_CONB_0;
  wire tie_lo_T10Y85__R2_CONB_0;
  wire tie_lo_T10Y86__R2_CONB_0;
  wire tie_lo_T10Y87__R2_CONB_0;
  wire tie_lo_T10Y88__R2_CONB_0;
  wire tie_lo_T10Y89__R2_CONB_0;
  wire tie_lo_T10Y8__R2_CONB_0;
  wire tie_lo_T10Y9__R2_CONB_0;
  wire tie_lo_T11Y0__R2_CONB_0;
  wire tie_lo_T11Y10__R2_CONB_0;
  wire tie_lo_T11Y11__R2_CONB_0;
  wire tie_lo_T11Y12__R2_CONB_0;
  wire tie_lo_T11Y13__R2_CONB_0;
  wire tie_lo_T11Y14__R2_CONB_0;
  wire tie_lo_T11Y15__R2_CONB_0;
  wire tie_lo_T11Y16__R2_CONB_0;
  wire tie_lo_T11Y17__R2_CONB_0;
  wire tie_lo_T11Y18__R2_CONB_0;
  wire tie_lo_T11Y19__R2_CONB_0;
  wire tie_lo_T11Y1__R2_CONB_0;
  wire tie_lo_T11Y20__R2_CONB_0;
  wire tie_lo_T11Y21__R2_CONB_0;
  wire tie_lo_T11Y22__R2_CONB_0;
  wire tie_lo_T11Y23__R2_CONB_0;
  wire tie_lo_T11Y24__R2_CONB_0;
  wire tie_lo_T11Y25__R2_CONB_0;
  wire tie_lo_T11Y26__R2_CONB_0;
  wire tie_lo_T11Y27__R2_CONB_0;
  wire tie_lo_T11Y28__R2_CONB_0;
  wire tie_lo_T11Y29__R2_CONB_0;
  wire tie_lo_T11Y2__R2_CONB_0;
  wire tie_lo_T11Y30__R2_CONB_0;
  wire tie_lo_T11Y31__R2_CONB_0;
  wire tie_lo_T11Y32__R2_CONB_0;
  wire tie_lo_T11Y33__R2_CONB_0;
  wire tie_lo_T11Y34__R2_CONB_0;
  wire tie_lo_T11Y35__R2_CONB_0;
  wire tie_lo_T11Y36__R2_CONB_0;
  wire tie_lo_T11Y37__R2_CONB_0;
  wire tie_lo_T11Y38__R2_CONB_0;
  wire tie_lo_T11Y39__R2_CONB_0;
  wire tie_lo_T11Y3__R2_CONB_0;
  wire tie_lo_T11Y40__R2_CONB_0;
  wire tie_lo_T11Y41__R2_CONB_0;
  wire tie_lo_T11Y42__R2_CONB_0;
  wire tie_lo_T11Y43__R2_CONB_0;
  wire tie_lo_T11Y44__R2_CONB_0;
  wire tie_lo_T11Y45__R2_CONB_0;
  wire tie_lo_T11Y46__R2_CONB_0;
  wire tie_lo_T11Y47__R2_CONB_0;
  wire tie_lo_T11Y48__R2_CONB_0;
  wire tie_lo_T11Y49__R2_CONB_0;
  wire tie_lo_T11Y4__R2_CONB_0;
  wire tie_lo_T11Y50__R2_CONB_0;
  wire tie_lo_T11Y51__R2_CONB_0;
  wire tie_lo_T11Y52__R2_CONB_0;
  wire tie_lo_T11Y53__R2_CONB_0;
  wire tie_lo_T11Y54__R2_CONB_0;
  wire tie_lo_T11Y55__R2_CONB_0;
  wire tie_lo_T11Y56__R2_CONB_0;
  wire tie_lo_T11Y57__R2_CONB_0;
  wire tie_lo_T11Y58__R2_CONB_0;
  wire tie_lo_T11Y59__R2_CONB_0;
  wire tie_lo_T11Y5__R2_CONB_0;
  wire tie_lo_T11Y60__R2_CONB_0;
  wire tie_lo_T11Y61__R2_CONB_0;
  wire tie_lo_T11Y62__R2_CONB_0;
  wire tie_lo_T11Y63__R2_CONB_0;
  wire tie_lo_T11Y64__R2_CONB_0;
  wire tie_lo_T11Y65__R2_CONB_0;
  wire tie_lo_T11Y66__R2_CONB_0;
  wire tie_lo_T11Y67__R2_CONB_0;
  wire tie_lo_T11Y68__R2_CONB_0;
  wire tie_lo_T11Y69__R2_CONB_0;
  wire tie_lo_T11Y6__R2_CONB_0;
  wire tie_lo_T11Y70__R2_CONB_0;
  wire tie_lo_T11Y71__R2_CONB_0;
  wire tie_lo_T11Y72__R2_CONB_0;
  wire tie_lo_T11Y73__R2_CONB_0;
  wire tie_lo_T11Y74__R2_CONB_0;
  wire tie_lo_T11Y75__R2_CONB_0;
  wire tie_lo_T11Y76__R2_CONB_0;
  wire tie_lo_T11Y77__R2_CONB_0;
  wire tie_lo_T11Y78__R2_CONB_0;
  wire tie_lo_T11Y79__R2_CONB_0;
  wire tie_lo_T11Y7__R2_CONB_0;
  wire tie_lo_T11Y80__R2_CONB_0;
  wire tie_lo_T11Y81__R2_CONB_0;
  wire tie_lo_T11Y82__R2_CONB_0;
  wire tie_lo_T11Y83__R2_CONB_0;
  wire tie_lo_T11Y84__R2_CONB_0;
  wire tie_lo_T11Y85__R2_CONB_0;
  wire tie_lo_T11Y86__R2_CONB_0;
  wire tie_lo_T11Y87__R2_CONB_0;
  wire tie_lo_T11Y88__R2_CONB_0;
  wire tie_lo_T11Y89__R2_CONB_0;
  wire tie_lo_T11Y8__R2_CONB_0;
  wire tie_lo_T11Y9__R2_CONB_0;
  wire tie_lo_T12Y0__R2_CONB_0;
  wire tie_lo_T12Y10__R2_CONB_0;
  wire tie_lo_T12Y11__R2_CONB_0;
  wire tie_lo_T12Y12__R2_CONB_0;
  wire tie_lo_T12Y13__R2_CONB_0;
  wire tie_lo_T12Y14__R2_CONB_0;
  wire tie_lo_T12Y15__R2_CONB_0;
  wire tie_lo_T12Y16__R2_CONB_0;
  wire tie_lo_T12Y17__R2_CONB_0;
  wire tie_lo_T12Y18__R2_CONB_0;
  wire tie_lo_T12Y19__R2_CONB_0;
  wire tie_lo_T12Y1__R2_CONB_0;
  wire tie_lo_T12Y20__R2_CONB_0;
  wire tie_lo_T12Y21__R2_CONB_0;
  wire tie_lo_T12Y22__R2_CONB_0;
  wire tie_lo_T12Y23__R2_CONB_0;
  wire tie_lo_T12Y24__R2_CONB_0;
  wire tie_lo_T12Y25__R2_CONB_0;
  wire tie_lo_T12Y26__R2_CONB_0;
  wire tie_lo_T12Y27__R2_CONB_0;
  wire tie_lo_T12Y28__R2_CONB_0;
  wire tie_lo_T12Y29__R2_CONB_0;
  wire tie_lo_T12Y2__R2_CONB_0;
  wire tie_lo_T12Y30__R2_CONB_0;
  wire tie_lo_T12Y31__R2_CONB_0;
  wire tie_lo_T12Y32__R2_CONB_0;
  wire tie_lo_T12Y33__R2_CONB_0;
  wire tie_lo_T12Y34__R2_CONB_0;
  wire tie_lo_T12Y35__R2_CONB_0;
  wire tie_lo_T12Y36__R2_CONB_0;
  wire tie_lo_T12Y37__R2_CONB_0;
  wire tie_lo_T12Y38__R2_CONB_0;
  wire tie_lo_T12Y39__R2_CONB_0;
  wire tie_lo_T12Y3__R2_CONB_0;
  wire tie_lo_T12Y40__R2_CONB_0;
  wire tie_lo_T12Y41__R2_CONB_0;
  wire tie_lo_T12Y42__R2_CONB_0;
  wire tie_lo_T12Y43__R2_CONB_0;
  wire tie_lo_T12Y44__R2_CONB_0;
  wire tie_lo_T12Y45__R2_CONB_0;
  wire tie_lo_T12Y46__R2_CONB_0;
  wire tie_lo_T12Y47__R2_CONB_0;
  wire tie_lo_T12Y48__R2_CONB_0;
  wire tie_lo_T12Y49__R2_CONB_0;
  wire tie_lo_T12Y4__R2_CONB_0;
  wire tie_lo_T12Y50__R2_CONB_0;
  wire tie_lo_T12Y51__R2_CONB_0;
  wire tie_lo_T12Y52__R2_CONB_0;
  wire tie_lo_T12Y53__R2_CONB_0;
  wire tie_lo_T12Y54__R2_CONB_0;
  wire tie_lo_T12Y55__R2_CONB_0;
  wire tie_lo_T12Y56__R2_CONB_0;
  wire tie_lo_T12Y57__R2_CONB_0;
  wire tie_lo_T12Y58__R2_CONB_0;
  wire tie_lo_T12Y59__R2_CONB_0;
  wire tie_lo_T12Y5__R2_CONB_0;
  wire tie_lo_T12Y60__R2_CONB_0;
  wire tie_lo_T12Y61__R2_CONB_0;
  wire tie_lo_T12Y62__R2_CONB_0;
  wire tie_lo_T12Y63__R2_CONB_0;
  wire tie_lo_T12Y64__R2_CONB_0;
  wire tie_lo_T12Y65__R2_CONB_0;
  wire tie_lo_T12Y66__R2_CONB_0;
  wire tie_lo_T12Y67__R2_CONB_0;
  wire tie_lo_T12Y68__R2_CONB_0;
  wire tie_lo_T12Y69__R2_CONB_0;
  wire tie_lo_T12Y6__R2_CONB_0;
  wire tie_lo_T12Y70__R2_CONB_0;
  wire tie_lo_T12Y71__R2_CONB_0;
  wire tie_lo_T12Y72__R2_CONB_0;
  wire tie_lo_T12Y73__R2_CONB_0;
  wire tie_lo_T12Y74__R2_CONB_0;
  wire tie_lo_T12Y75__R2_CONB_0;
  wire tie_lo_T12Y76__R2_CONB_0;
  wire tie_lo_T12Y77__R2_CONB_0;
  wire tie_lo_T12Y78__R2_CONB_0;
  wire tie_lo_T12Y79__R2_CONB_0;
  wire tie_lo_T12Y7__R2_CONB_0;
  wire tie_lo_T12Y80__R2_CONB_0;
  wire tie_lo_T12Y81__R2_CONB_0;
  wire tie_lo_T12Y82__R2_CONB_0;
  wire tie_lo_T12Y83__R2_CONB_0;
  wire tie_lo_T12Y84__R2_CONB_0;
  wire tie_lo_T12Y85__R2_CONB_0;
  wire tie_lo_T12Y86__R2_CONB_0;
  wire tie_lo_T12Y87__R2_CONB_0;
  wire tie_lo_T12Y88__R2_CONB_0;
  wire tie_lo_T12Y89__R2_CONB_0;
  wire tie_lo_T12Y8__R2_CONB_0;
  wire tie_lo_T12Y9__R2_CONB_0;
  wire tie_lo_T13Y0__R2_CONB_0;
  wire tie_lo_T13Y10__R2_CONB_0;
  wire tie_lo_T13Y11__R2_CONB_0;
  wire tie_lo_T13Y12__R2_CONB_0;
  wire tie_lo_T13Y13__R2_CONB_0;
  wire tie_lo_T13Y14__R2_CONB_0;
  wire tie_lo_T13Y15__R2_CONB_0;
  wire tie_lo_T13Y16__R2_CONB_0;
  wire tie_lo_T13Y17__R2_CONB_0;
  wire tie_lo_T13Y18__R2_CONB_0;
  wire tie_lo_T13Y19__R2_CONB_0;
  wire tie_lo_T13Y1__R2_CONB_0;
  wire tie_lo_T13Y20__R2_CONB_0;
  wire tie_lo_T13Y21__R2_CONB_0;
  wire tie_lo_T13Y22__R2_CONB_0;
  wire tie_lo_T13Y23__R2_CONB_0;
  wire tie_lo_T13Y24__R2_CONB_0;
  wire tie_lo_T13Y25__R2_CONB_0;
  wire tie_lo_T13Y26__R2_CONB_0;
  wire tie_lo_T13Y27__R2_CONB_0;
  wire tie_lo_T13Y28__R2_CONB_0;
  wire tie_lo_T13Y29__R2_CONB_0;
  wire tie_lo_T13Y2__R2_CONB_0;
  wire tie_lo_T13Y30__R2_CONB_0;
  wire tie_lo_T13Y31__R2_CONB_0;
  wire tie_lo_T13Y32__R2_CONB_0;
  wire tie_lo_T13Y33__R2_CONB_0;
  wire tie_lo_T13Y34__R2_CONB_0;
  wire tie_lo_T13Y35__R2_CONB_0;
  wire tie_lo_T13Y36__R2_CONB_0;
  wire tie_lo_T13Y37__R2_CONB_0;
  wire tie_lo_T13Y38__R2_CONB_0;
  wire tie_lo_T13Y39__R2_CONB_0;
  wire tie_lo_T13Y3__R2_CONB_0;
  wire tie_lo_T13Y40__R2_CONB_0;
  wire tie_lo_T13Y41__R2_CONB_0;
  wire tie_lo_T13Y42__R2_CONB_0;
  wire tie_lo_T13Y43__R2_CONB_0;
  wire tie_lo_T13Y44__R2_CONB_0;
  wire tie_lo_T13Y45__R2_CONB_0;
  wire tie_lo_T13Y46__R2_CONB_0;
  wire tie_lo_T13Y47__R2_CONB_0;
  wire tie_lo_T13Y48__R2_CONB_0;
  wire tie_lo_T13Y49__R2_CONB_0;
  wire tie_lo_T13Y4__R2_CONB_0;
  wire tie_lo_T13Y50__R2_CONB_0;
  wire tie_lo_T13Y51__R2_CONB_0;
  wire tie_lo_T13Y52__R2_CONB_0;
  wire tie_lo_T13Y53__R2_CONB_0;
  wire tie_lo_T13Y54__R2_CONB_0;
  wire tie_lo_T13Y55__R2_CONB_0;
  wire tie_lo_T13Y56__R2_CONB_0;
  wire tie_lo_T13Y57__R2_CONB_0;
  wire tie_lo_T13Y58__R2_CONB_0;
  wire tie_lo_T13Y59__R2_CONB_0;
  wire tie_lo_T13Y5__R2_CONB_0;
  wire tie_lo_T13Y60__R2_CONB_0;
  wire tie_lo_T13Y61__R2_CONB_0;
  wire tie_lo_T13Y62__R2_CONB_0;
  wire tie_lo_T13Y63__R2_CONB_0;
  wire tie_lo_T13Y64__R2_CONB_0;
  wire tie_lo_T13Y65__R2_CONB_0;
  wire tie_lo_T13Y66__R2_CONB_0;
  wire tie_lo_T13Y67__R2_CONB_0;
  wire tie_lo_T13Y68__R2_CONB_0;
  wire tie_lo_T13Y69__R2_CONB_0;
  wire tie_lo_T13Y6__R2_CONB_0;
  wire tie_lo_T13Y70__R2_CONB_0;
  wire tie_lo_T13Y71__R2_CONB_0;
  wire tie_lo_T13Y72__R2_CONB_0;
  wire tie_lo_T13Y73__R2_CONB_0;
  wire tie_lo_T13Y74__R2_CONB_0;
  wire tie_lo_T13Y75__R2_CONB_0;
  wire tie_lo_T13Y76__R2_CONB_0;
  wire tie_lo_T13Y77__R2_CONB_0;
  wire tie_lo_T13Y78__R2_CONB_0;
  wire tie_lo_T13Y79__R2_CONB_0;
  wire tie_lo_T13Y7__R2_CONB_0;
  wire tie_lo_T13Y80__R2_CONB_0;
  wire tie_lo_T13Y81__R2_CONB_0;
  wire tie_lo_T13Y82__R2_CONB_0;
  wire tie_lo_T13Y83__R2_CONB_0;
  wire tie_lo_T13Y84__R2_CONB_0;
  wire tie_lo_T13Y85__R2_CONB_0;
  wire tie_lo_T13Y86__R2_CONB_0;
  wire tie_lo_T13Y87__R2_CONB_0;
  wire tie_lo_T13Y88__R2_CONB_0;
  wire tie_lo_T13Y89__R2_CONB_0;
  wire tie_lo_T13Y8__R2_CONB_0;
  wire tie_lo_T13Y9__R2_CONB_0;
  wire tie_lo_T14Y0__R2_CONB_0;
  wire tie_lo_T14Y10__R2_CONB_0;
  wire tie_lo_T14Y11__R2_CONB_0;
  wire tie_lo_T14Y12__R2_CONB_0;
  wire tie_lo_T14Y13__R2_CONB_0;
  wire tie_lo_T14Y14__R2_CONB_0;
  wire tie_lo_T14Y15__R2_CONB_0;
  wire tie_lo_T14Y16__R2_CONB_0;
  wire tie_lo_T14Y17__R2_CONB_0;
  wire tie_lo_T14Y18__R2_CONB_0;
  wire tie_lo_T14Y19__R2_CONB_0;
  wire tie_lo_T14Y1__R2_CONB_0;
  wire tie_lo_T14Y20__R2_CONB_0;
  wire tie_lo_T14Y21__R2_CONB_0;
  wire tie_lo_T14Y22__R2_CONB_0;
  wire tie_lo_T14Y23__R2_CONB_0;
  wire tie_lo_T14Y24__R2_CONB_0;
  wire tie_lo_T14Y25__R2_CONB_0;
  wire tie_lo_T14Y26__R2_CONB_0;
  wire tie_lo_T14Y27__R2_CONB_0;
  wire tie_lo_T14Y28__R2_CONB_0;
  wire tie_lo_T14Y29__R2_CONB_0;
  wire tie_lo_T14Y2__R2_CONB_0;
  wire tie_lo_T14Y30__R2_CONB_0;
  wire tie_lo_T14Y31__R2_CONB_0;
  wire tie_lo_T14Y32__R2_CONB_0;
  wire tie_lo_T14Y33__R2_CONB_0;
  wire tie_lo_T14Y34__R2_CONB_0;
  wire tie_lo_T14Y35__R2_CONB_0;
  wire tie_lo_T14Y36__R2_CONB_0;
  wire tie_lo_T14Y37__R2_CONB_0;
  wire tie_lo_T14Y38__R2_CONB_0;
  wire tie_lo_T14Y39__R2_CONB_0;
  wire tie_lo_T14Y3__R2_CONB_0;
  wire tie_lo_T14Y40__R2_CONB_0;
  wire tie_lo_T14Y41__R2_CONB_0;
  wire tie_lo_T14Y42__R2_CONB_0;
  wire tie_lo_T14Y43__R2_CONB_0;
  wire tie_lo_T14Y44__R2_CONB_0;
  wire tie_lo_T14Y45__R2_CONB_0;
  wire tie_lo_T14Y46__R2_CONB_0;
  wire tie_lo_T14Y47__R2_CONB_0;
  wire tie_lo_T14Y48__R2_CONB_0;
  wire tie_lo_T14Y49__R2_CONB_0;
  wire tie_lo_T14Y4__R2_CONB_0;
  wire tie_lo_T14Y50__R2_CONB_0;
  wire tie_lo_T14Y51__R2_CONB_0;
  wire tie_lo_T14Y52__R2_CONB_0;
  wire tie_lo_T14Y53__R2_CONB_0;
  wire tie_lo_T14Y54__R2_CONB_0;
  wire tie_lo_T14Y55__R2_CONB_0;
  wire tie_lo_T14Y56__R2_CONB_0;
  wire tie_lo_T14Y57__R2_CONB_0;
  wire tie_lo_T14Y58__R2_CONB_0;
  wire tie_lo_T14Y59__R2_CONB_0;
  wire tie_lo_T14Y5__R2_CONB_0;
  wire tie_lo_T14Y60__R2_CONB_0;
  wire tie_lo_T14Y61__R2_CONB_0;
  wire tie_lo_T14Y62__R2_CONB_0;
  wire tie_lo_T14Y63__R2_CONB_0;
  wire tie_lo_T14Y64__R2_CONB_0;
  wire tie_lo_T14Y65__R2_CONB_0;
  wire tie_lo_T14Y66__R2_CONB_0;
  wire tie_lo_T14Y67__R2_CONB_0;
  wire tie_lo_T14Y68__R2_CONB_0;
  wire tie_lo_T14Y69__R2_CONB_0;
  wire tie_lo_T14Y6__R2_CONB_0;
  wire tie_lo_T14Y70__R2_CONB_0;
  wire tie_lo_T14Y71__R2_CONB_0;
  wire tie_lo_T14Y72__R2_CONB_0;
  wire tie_lo_T14Y73__R2_CONB_0;
  wire tie_lo_T14Y74__R2_CONB_0;
  wire tie_lo_T14Y75__R2_CONB_0;
  wire tie_lo_T14Y76__R2_CONB_0;
  wire tie_lo_T14Y77__R2_CONB_0;
  wire tie_lo_T14Y78__R2_CONB_0;
  wire tie_lo_T14Y79__R2_CONB_0;
  wire tie_lo_T14Y7__R2_CONB_0;
  wire tie_lo_T14Y80__R2_CONB_0;
  wire tie_lo_T14Y81__R2_CONB_0;
  wire tie_lo_T14Y82__R2_CONB_0;
  wire tie_lo_T14Y83__R2_CONB_0;
  wire tie_lo_T14Y84__R2_CONB_0;
  wire tie_lo_T14Y85__R2_CONB_0;
  wire tie_lo_T14Y86__R2_CONB_0;
  wire tie_lo_T14Y87__R2_CONB_0;
  wire tie_lo_T14Y88__R2_CONB_0;
  wire tie_lo_T14Y89__R2_CONB_0;
  wire tie_lo_T14Y8__R2_CONB_0;
  wire tie_lo_T14Y9__R2_CONB_0;
  wire tie_lo_T15Y0__R2_CONB_0;
  wire tie_lo_T15Y10__R2_CONB_0;
  wire tie_lo_T15Y11__R2_CONB_0;
  wire tie_lo_T15Y12__R2_CONB_0;
  wire tie_lo_T15Y13__R2_CONB_0;
  wire tie_lo_T15Y14__R2_CONB_0;
  wire tie_lo_T15Y15__R2_CONB_0;
  wire tie_lo_T15Y16__R2_CONB_0;
  wire tie_lo_T15Y17__R2_CONB_0;
  wire tie_lo_T15Y18__R2_CONB_0;
  wire tie_lo_T15Y19__R2_CONB_0;
  wire tie_lo_T15Y1__R2_CONB_0;
  wire tie_lo_T15Y20__R2_CONB_0;
  wire tie_lo_T15Y21__R2_CONB_0;
  wire tie_lo_T15Y22__R2_CONB_0;
  wire tie_lo_T15Y23__R2_CONB_0;
  wire tie_lo_T15Y24__R2_CONB_0;
  wire tie_lo_T15Y25__R2_CONB_0;
  wire tie_lo_T15Y26__R2_CONB_0;
  wire tie_lo_T15Y27__R2_CONB_0;
  wire tie_lo_T15Y28__R2_CONB_0;
  wire tie_lo_T15Y29__R2_CONB_0;
  wire tie_lo_T15Y2__R2_CONB_0;
  wire tie_lo_T15Y30__R2_CONB_0;
  wire tie_lo_T15Y31__R2_CONB_0;
  wire tie_lo_T15Y32__R2_CONB_0;
  wire tie_lo_T15Y33__R2_CONB_0;
  wire tie_lo_T15Y34__R2_CONB_0;
  wire tie_lo_T15Y35__R2_CONB_0;
  wire tie_lo_T15Y36__R2_CONB_0;
  wire tie_lo_T15Y37__R2_CONB_0;
  wire tie_lo_T15Y38__R2_CONB_0;
  wire tie_lo_T15Y39__R2_CONB_0;
  wire tie_lo_T15Y3__R2_CONB_0;
  wire tie_lo_T15Y40__R2_CONB_0;
  wire tie_lo_T15Y41__R2_CONB_0;
  wire tie_lo_T15Y42__R2_CONB_0;
  wire tie_lo_T15Y43__R2_CONB_0;
  wire tie_lo_T15Y44__R2_CONB_0;
  wire tie_lo_T15Y45__R2_CONB_0;
  wire tie_lo_T15Y46__R2_CONB_0;
  wire tie_lo_T15Y47__R2_CONB_0;
  wire tie_lo_T15Y48__R2_CONB_0;
  wire tie_lo_T15Y49__R2_CONB_0;
  wire tie_lo_T15Y4__R2_CONB_0;
  wire tie_lo_T15Y50__R2_CONB_0;
  wire tie_lo_T15Y51__R2_CONB_0;
  wire tie_lo_T15Y52__R2_CONB_0;
  wire tie_lo_T15Y53__R2_CONB_0;
  wire tie_lo_T15Y54__R2_CONB_0;
  wire tie_lo_T15Y55__R2_CONB_0;
  wire tie_lo_T15Y56__R2_CONB_0;
  wire tie_lo_T15Y57__R2_CONB_0;
  wire tie_lo_T15Y58__R2_CONB_0;
  wire tie_lo_T15Y59__R2_CONB_0;
  wire tie_lo_T15Y5__R2_CONB_0;
  wire tie_lo_T15Y60__R2_CONB_0;
  wire tie_lo_T15Y61__R2_CONB_0;
  wire tie_lo_T15Y62__R2_CONB_0;
  wire tie_lo_T15Y63__R2_CONB_0;
  wire tie_lo_T15Y64__R2_CONB_0;
  wire tie_lo_T15Y65__R2_CONB_0;
  wire tie_lo_T15Y66__R2_CONB_0;
  wire tie_lo_T15Y67__R2_CONB_0;
  wire tie_lo_T15Y68__R2_CONB_0;
  wire tie_lo_T15Y69__R2_CONB_0;
  wire tie_lo_T15Y6__R2_CONB_0;
  wire tie_lo_T15Y70__R2_CONB_0;
  wire tie_lo_T15Y71__R2_CONB_0;
  wire tie_lo_T15Y72__R2_CONB_0;
  wire tie_lo_T15Y73__R2_CONB_0;
  wire tie_lo_T15Y74__R2_CONB_0;
  wire tie_lo_T15Y75__R2_CONB_0;
  wire tie_lo_T15Y76__R2_CONB_0;
  wire tie_lo_T15Y77__R2_CONB_0;
  wire tie_lo_T15Y78__R2_CONB_0;
  wire tie_lo_T15Y79__R2_CONB_0;
  wire tie_lo_T15Y7__R2_CONB_0;
  wire tie_lo_T15Y80__R2_CONB_0;
  wire tie_lo_T15Y81__R2_CONB_0;
  wire tie_lo_T15Y82__R2_CONB_0;
  wire tie_lo_T15Y83__R2_CONB_0;
  wire tie_lo_T15Y84__R2_CONB_0;
  wire tie_lo_T15Y85__R2_CONB_0;
  wire tie_lo_T15Y86__R2_CONB_0;
  wire tie_lo_T15Y87__R2_CONB_0;
  wire tie_lo_T15Y88__R2_CONB_0;
  wire tie_lo_T15Y89__R2_CONB_0;
  wire tie_lo_T15Y8__R2_CONB_0;
  wire tie_lo_T15Y9__R2_CONB_0;
  wire tie_lo_T16Y0__R2_CONB_0;
  wire tie_lo_T16Y10__R2_CONB_0;
  wire tie_lo_T16Y11__R2_CONB_0;
  wire tie_lo_T16Y12__R2_CONB_0;
  wire tie_lo_T16Y13__R2_CONB_0;
  wire tie_lo_T16Y14__R2_CONB_0;
  wire tie_lo_T16Y15__R2_CONB_0;
  wire tie_lo_T16Y16__R2_CONB_0;
  wire tie_lo_T16Y17__R2_CONB_0;
  wire tie_lo_T16Y18__R2_CONB_0;
  wire tie_lo_T16Y19__R2_CONB_0;
  wire tie_lo_T16Y1__R2_CONB_0;
  wire tie_lo_T16Y20__R2_CONB_0;
  wire tie_lo_T16Y21__R2_CONB_0;
  wire tie_lo_T16Y22__R2_CONB_0;
  wire tie_lo_T16Y23__R2_CONB_0;
  wire tie_lo_T16Y24__R2_CONB_0;
  wire tie_lo_T16Y25__R2_CONB_0;
  wire tie_lo_T16Y26__R2_CONB_0;
  wire tie_lo_T16Y27__R2_CONB_0;
  wire tie_lo_T16Y28__R2_CONB_0;
  wire tie_lo_T16Y29__R2_CONB_0;
  wire tie_lo_T16Y2__R2_CONB_0;
  wire tie_lo_T16Y30__R2_CONB_0;
  wire tie_lo_T16Y31__R2_CONB_0;
  wire tie_lo_T16Y32__R2_CONB_0;
  wire tie_lo_T16Y33__R2_CONB_0;
  wire tie_lo_T16Y34__R2_CONB_0;
  wire tie_lo_T16Y35__R2_CONB_0;
  wire tie_lo_T16Y36__R2_CONB_0;
  wire tie_lo_T16Y37__R2_CONB_0;
  wire tie_lo_T16Y38__R2_CONB_0;
  wire tie_lo_T16Y39__R2_CONB_0;
  wire tie_lo_T16Y3__R2_CONB_0;
  wire tie_lo_T16Y40__R2_CONB_0;
  wire tie_lo_T16Y41__R2_CONB_0;
  wire tie_lo_T16Y42__R2_CONB_0;
  wire tie_lo_T16Y43__R2_CONB_0;
  wire tie_lo_T16Y44__R2_CONB_0;
  wire tie_lo_T16Y45__R2_CONB_0;
  wire tie_lo_T16Y46__R2_CONB_0;
  wire tie_lo_T16Y47__R2_CONB_0;
  wire tie_lo_T16Y48__R2_CONB_0;
  wire tie_lo_T16Y49__R2_CONB_0;
  wire tie_lo_T16Y4__R2_CONB_0;
  wire tie_lo_T16Y50__R2_CONB_0;
  wire tie_lo_T16Y51__R2_CONB_0;
  wire tie_lo_T16Y52__R2_CONB_0;
  wire tie_lo_T16Y53__R2_CONB_0;
  wire tie_lo_T16Y54__R2_CONB_0;
  wire tie_lo_T16Y55__R2_CONB_0;
  wire tie_lo_T16Y56__R2_CONB_0;
  wire tie_lo_T16Y57__R2_CONB_0;
  wire tie_lo_T16Y58__R2_CONB_0;
  wire tie_lo_T16Y59__R2_CONB_0;
  wire tie_lo_T16Y5__R2_CONB_0;
  wire tie_lo_T16Y60__R2_CONB_0;
  wire tie_lo_T16Y61__R2_CONB_0;
  wire tie_lo_T16Y62__R2_CONB_0;
  wire tie_lo_T16Y63__R2_CONB_0;
  wire tie_lo_T16Y64__R2_CONB_0;
  wire tie_lo_T16Y65__R2_CONB_0;
  wire tie_lo_T16Y66__R2_CONB_0;
  wire tie_lo_T16Y67__R2_CONB_0;
  wire tie_lo_T16Y68__R2_CONB_0;
  wire tie_lo_T16Y69__R2_CONB_0;
  wire tie_lo_T16Y6__R2_CONB_0;
  wire tie_lo_T16Y70__R2_CONB_0;
  wire tie_lo_T16Y71__R2_CONB_0;
  wire tie_lo_T16Y72__R2_CONB_0;
  wire tie_lo_T16Y73__R2_CONB_0;
  wire tie_lo_T16Y74__R2_CONB_0;
  wire tie_lo_T16Y75__R2_CONB_0;
  wire tie_lo_T16Y76__R2_CONB_0;
  wire tie_lo_T16Y77__R2_CONB_0;
  wire tie_lo_T16Y78__R2_CONB_0;
  wire tie_lo_T16Y79__R2_CONB_0;
  wire tie_lo_T16Y7__R2_CONB_0;
  wire tie_lo_T16Y80__R2_CONB_0;
  wire tie_lo_T16Y81__R2_CONB_0;
  wire tie_lo_T16Y82__R2_CONB_0;
  wire tie_lo_T16Y83__R2_CONB_0;
  wire tie_lo_T16Y84__R2_CONB_0;
  wire tie_lo_T16Y85__R2_CONB_0;
  wire tie_lo_T16Y86__R2_CONB_0;
  wire tie_lo_T16Y87__R2_CONB_0;
  wire tie_lo_T16Y88__R2_CONB_0;
  wire tie_lo_T16Y89__R2_CONB_0;
  wire tie_lo_T16Y8__R2_CONB_0;
  wire tie_lo_T16Y9__R2_CONB_0;
  wire tie_lo_T17Y0__R2_CONB_0;
  wire tie_lo_T17Y10__R2_CONB_0;
  wire tie_lo_T17Y11__R2_CONB_0;
  wire tie_lo_T17Y12__R2_CONB_0;
  wire tie_lo_T17Y13__R2_CONB_0;
  wire tie_lo_T17Y14__R2_CONB_0;
  wire tie_lo_T17Y15__R2_CONB_0;
  wire tie_lo_T17Y16__R2_CONB_0;
  wire tie_lo_T17Y17__R2_CONB_0;
  wire tie_lo_T17Y18__R2_CONB_0;
  wire tie_lo_T17Y19__R2_CONB_0;
  wire tie_lo_T17Y1__R2_CONB_0;
  wire tie_lo_T17Y20__R2_CONB_0;
  wire tie_lo_T17Y21__R2_CONB_0;
  wire tie_lo_T17Y22__R2_CONB_0;
  wire tie_lo_T17Y23__R2_CONB_0;
  wire tie_lo_T17Y24__R2_CONB_0;
  wire tie_lo_T17Y25__R2_CONB_0;
  wire tie_lo_T17Y26__R2_CONB_0;
  wire tie_lo_T17Y27__R2_CONB_0;
  wire tie_lo_T17Y28__R2_CONB_0;
  wire tie_lo_T17Y29__R2_CONB_0;
  wire tie_lo_T17Y2__R2_CONB_0;
  wire tie_lo_T17Y30__R2_CONB_0;
  wire tie_lo_T17Y31__R2_CONB_0;
  wire tie_lo_T17Y32__R2_CONB_0;
  wire tie_lo_T17Y33__R2_CONB_0;
  wire tie_lo_T17Y34__R2_CONB_0;
  wire tie_lo_T17Y35__R2_CONB_0;
  wire tie_lo_T17Y36__R2_CONB_0;
  wire tie_lo_T17Y37__R2_CONB_0;
  wire tie_lo_T17Y38__R2_CONB_0;
  wire tie_lo_T17Y39__R2_CONB_0;
  wire tie_lo_T17Y3__R2_CONB_0;
  wire tie_lo_T17Y40__R2_CONB_0;
  wire tie_lo_T17Y41__R2_CONB_0;
  wire tie_lo_T17Y42__R2_CONB_0;
  wire tie_lo_T17Y43__R2_CONB_0;
  wire tie_lo_T17Y44__R2_CONB_0;
  wire tie_lo_T17Y45__R2_CONB_0;
  wire tie_lo_T17Y46__R2_CONB_0;
  wire tie_lo_T17Y47__R2_CONB_0;
  wire tie_lo_T17Y48__R2_CONB_0;
  wire tie_lo_T17Y49__R2_CONB_0;
  wire tie_lo_T17Y4__R2_CONB_0;
  wire tie_lo_T17Y50__R2_CONB_0;
  wire tie_lo_T17Y51__R2_CONB_0;
  wire tie_lo_T17Y52__R2_CONB_0;
  wire tie_lo_T17Y53__R2_CONB_0;
  wire tie_lo_T17Y54__R2_CONB_0;
  wire tie_lo_T17Y55__R2_CONB_0;
  wire tie_lo_T17Y56__R2_CONB_0;
  wire tie_lo_T17Y57__R2_CONB_0;
  wire tie_lo_T17Y58__R2_CONB_0;
  wire tie_lo_T17Y59__R2_CONB_0;
  wire tie_lo_T17Y5__R2_CONB_0;
  wire tie_lo_T17Y60__R2_CONB_0;
  wire tie_lo_T17Y61__R2_CONB_0;
  wire tie_lo_T17Y62__R2_CONB_0;
  wire tie_lo_T17Y63__R2_CONB_0;
  wire tie_lo_T17Y64__R2_CONB_0;
  wire tie_lo_T17Y65__R2_CONB_0;
  wire tie_lo_T17Y66__R2_CONB_0;
  wire tie_lo_T17Y67__R2_CONB_0;
  wire tie_lo_T17Y68__R2_CONB_0;
  wire tie_lo_T17Y69__R2_CONB_0;
  wire tie_lo_T17Y6__R2_CONB_0;
  wire tie_lo_T17Y70__R2_CONB_0;
  wire tie_lo_T17Y71__R2_CONB_0;
  wire tie_lo_T17Y72__R2_CONB_0;
  wire tie_lo_T17Y73__R2_CONB_0;
  wire tie_lo_T17Y74__R2_CONB_0;
  wire tie_lo_T17Y75__R2_CONB_0;
  wire tie_lo_T17Y76__R2_CONB_0;
  wire tie_lo_T17Y77__R2_CONB_0;
  wire tie_lo_T17Y78__R2_CONB_0;
  wire tie_lo_T17Y79__R2_CONB_0;
  wire tie_lo_T17Y7__R2_CONB_0;
  wire tie_lo_T17Y80__R2_CONB_0;
  wire tie_lo_T17Y81__R2_CONB_0;
  wire tie_lo_T17Y82__R2_CONB_0;
  wire tie_lo_T17Y83__R2_CONB_0;
  wire tie_lo_T17Y84__R2_CONB_0;
  wire tie_lo_T17Y85__R2_CONB_0;
  wire tie_lo_T17Y86__R2_CONB_0;
  wire tie_lo_T17Y87__R2_CONB_0;
  wire tie_lo_T17Y88__R2_CONB_0;
  wire tie_lo_T17Y89__R2_CONB_0;
  wire tie_lo_T17Y8__R2_CONB_0;
  wire tie_lo_T17Y9__R2_CONB_0;
  wire tie_lo_T18Y0__R2_CONB_0;
  wire tie_lo_T18Y10__R2_CONB_0;
  wire tie_lo_T18Y11__R2_CONB_0;
  wire tie_lo_T18Y12__R2_CONB_0;
  wire tie_lo_T18Y13__R2_CONB_0;
  wire tie_lo_T18Y14__R2_CONB_0;
  wire tie_lo_T18Y15__R2_CONB_0;
  wire tie_lo_T18Y16__R2_CONB_0;
  wire tie_lo_T18Y17__R2_CONB_0;
  wire tie_lo_T18Y18__R2_CONB_0;
  wire tie_lo_T18Y19__R2_CONB_0;
  wire tie_lo_T18Y1__R2_CONB_0;
  wire tie_lo_T18Y20__R2_CONB_0;
  wire tie_lo_T18Y21__R2_CONB_0;
  wire tie_lo_T18Y22__R2_CONB_0;
  wire tie_lo_T18Y23__R2_CONB_0;
  wire tie_lo_T18Y24__R2_CONB_0;
  wire tie_lo_T18Y25__R2_CONB_0;
  wire tie_lo_T18Y26__R2_CONB_0;
  wire tie_lo_T18Y27__R2_CONB_0;
  wire tie_lo_T18Y28__R2_CONB_0;
  wire tie_lo_T18Y29__R2_CONB_0;
  wire tie_lo_T18Y2__R2_CONB_0;
  wire tie_lo_T18Y30__R2_CONB_0;
  wire tie_lo_T18Y31__R2_CONB_0;
  wire tie_lo_T18Y32__R2_CONB_0;
  wire tie_lo_T18Y33__R2_CONB_0;
  wire tie_lo_T18Y34__R2_CONB_0;
  wire tie_lo_T18Y35__R2_CONB_0;
  wire tie_lo_T18Y36__R2_CONB_0;
  wire tie_lo_T18Y37__R2_CONB_0;
  wire tie_lo_T18Y38__R2_CONB_0;
  wire tie_lo_T18Y39__R2_CONB_0;
  wire tie_lo_T18Y3__R2_CONB_0;
  wire tie_lo_T18Y40__R2_CONB_0;
  wire tie_lo_T18Y41__R2_CONB_0;
  wire tie_lo_T18Y42__R2_CONB_0;
  wire tie_lo_T18Y43__R2_CONB_0;
  wire tie_lo_T18Y44__R2_CONB_0;
  wire tie_lo_T18Y45__R2_CONB_0;
  wire tie_lo_T18Y46__R2_CONB_0;
  wire tie_lo_T18Y47__R2_CONB_0;
  wire tie_lo_T18Y48__R2_CONB_0;
  wire tie_lo_T18Y49__R2_CONB_0;
  wire tie_lo_T18Y4__R2_CONB_0;
  wire tie_lo_T18Y50__R2_CONB_0;
  wire tie_lo_T18Y51__R2_CONB_0;
  wire tie_lo_T18Y52__R2_CONB_0;
  wire tie_lo_T18Y53__R2_CONB_0;
  wire tie_lo_T18Y54__R2_CONB_0;
  wire tie_lo_T18Y55__R2_CONB_0;
  wire tie_lo_T18Y56__R2_CONB_0;
  wire tie_lo_T18Y57__R2_CONB_0;
  wire tie_lo_T18Y58__R2_CONB_0;
  wire tie_lo_T18Y59__R2_CONB_0;
  wire tie_lo_T18Y5__R2_CONB_0;
  wire tie_lo_T18Y60__R2_CONB_0;
  wire tie_lo_T18Y61__R2_CONB_0;
  wire tie_lo_T18Y62__R2_CONB_0;
  wire tie_lo_T18Y63__R2_CONB_0;
  wire tie_lo_T18Y64__R2_CONB_0;
  wire tie_lo_T18Y65__R2_CONB_0;
  wire tie_lo_T18Y66__R2_CONB_0;
  wire tie_lo_T18Y67__R2_CONB_0;
  wire tie_lo_T18Y68__R2_CONB_0;
  wire tie_lo_T18Y69__R2_CONB_0;
  wire tie_lo_T18Y6__R2_CONB_0;
  wire tie_lo_T18Y70__R2_CONB_0;
  wire tie_lo_T18Y71__R2_CONB_0;
  wire tie_lo_T18Y72__R2_CONB_0;
  wire tie_lo_T18Y73__R2_CONB_0;
  wire tie_lo_T18Y74__R2_CONB_0;
  wire tie_lo_T18Y75__R2_CONB_0;
  wire tie_lo_T18Y76__R2_CONB_0;
  wire tie_lo_T18Y77__R2_CONB_0;
  wire tie_lo_T18Y78__R2_CONB_0;
  wire tie_lo_T18Y79__R2_CONB_0;
  wire tie_lo_T18Y7__R2_CONB_0;
  wire tie_lo_T18Y80__R2_CONB_0;
  wire tie_lo_T18Y81__R2_CONB_0;
  wire tie_lo_T18Y82__R2_CONB_0;
  wire tie_lo_T18Y83__R2_CONB_0;
  wire tie_lo_T18Y84__R2_CONB_0;
  wire tie_lo_T18Y85__R2_CONB_0;
  wire tie_lo_T18Y86__R2_CONB_0;
  wire tie_lo_T18Y87__R2_CONB_0;
  wire tie_lo_T18Y88__R2_CONB_0;
  wire tie_lo_T18Y89__R2_CONB_0;
  wire tie_lo_T18Y8__R2_CONB_0;
  wire tie_lo_T18Y9__R2_CONB_0;
  wire tie_lo_T19Y0__R2_CONB_0;
  wire tie_lo_T19Y10__R2_CONB_0;
  wire tie_lo_T19Y11__R2_CONB_0;
  wire tie_lo_T19Y12__R2_CONB_0;
  wire tie_lo_T19Y13__R2_CONB_0;
  wire tie_lo_T19Y14__R2_CONB_0;
  wire tie_lo_T19Y15__R2_CONB_0;
  wire tie_lo_T19Y16__R2_CONB_0;
  wire tie_lo_T19Y17__R2_CONB_0;
  wire tie_lo_T19Y18__R2_CONB_0;
  wire tie_lo_T19Y19__R2_CONB_0;
  wire tie_lo_T19Y1__R2_CONB_0;
  wire tie_lo_T19Y20__R2_CONB_0;
  wire tie_lo_T19Y21__R2_CONB_0;
  wire tie_lo_T19Y22__R2_CONB_0;
  wire tie_lo_T19Y23__R2_CONB_0;
  wire tie_lo_T19Y24__R2_CONB_0;
  wire tie_lo_T19Y25__R2_CONB_0;
  wire tie_lo_T19Y26__R2_CONB_0;
  wire tie_lo_T19Y27__R2_CONB_0;
  wire tie_lo_T19Y28__R2_CONB_0;
  wire tie_lo_T19Y29__R2_CONB_0;
  wire tie_lo_T19Y2__R2_CONB_0;
  wire tie_lo_T19Y30__R2_CONB_0;
  wire tie_lo_T19Y31__R2_CONB_0;
  wire tie_lo_T19Y32__R2_CONB_0;
  wire tie_lo_T19Y33__R2_CONB_0;
  wire tie_lo_T19Y34__R2_CONB_0;
  wire tie_lo_T19Y35__R2_CONB_0;
  wire tie_lo_T19Y36__R2_CONB_0;
  wire tie_lo_T19Y37__R2_CONB_0;
  wire tie_lo_T19Y38__R2_CONB_0;
  wire tie_lo_T19Y39__R2_CONB_0;
  wire tie_lo_T19Y3__R2_CONB_0;
  wire tie_lo_T19Y40__R2_CONB_0;
  wire tie_lo_T19Y41__R2_CONB_0;
  wire tie_lo_T19Y42__R2_CONB_0;
  wire tie_lo_T19Y43__R2_CONB_0;
  wire tie_lo_T19Y44__R2_CONB_0;
  wire tie_lo_T19Y45__R2_CONB_0;
  wire tie_lo_T19Y46__R2_CONB_0;
  wire tie_lo_T19Y47__R2_CONB_0;
  wire tie_lo_T19Y48__R2_CONB_0;
  wire tie_lo_T19Y49__R2_CONB_0;
  wire tie_lo_T19Y4__R2_CONB_0;
  wire tie_lo_T19Y50__R2_CONB_0;
  wire tie_lo_T19Y51__R2_CONB_0;
  wire tie_lo_T19Y52__R2_CONB_0;
  wire tie_lo_T19Y53__R2_CONB_0;
  wire tie_lo_T19Y54__R2_CONB_0;
  wire tie_lo_T19Y55__R2_CONB_0;
  wire tie_lo_T19Y56__R2_CONB_0;
  wire tie_lo_T19Y57__R2_CONB_0;
  wire tie_lo_T19Y58__R2_CONB_0;
  wire tie_lo_T19Y59__R2_CONB_0;
  wire tie_lo_T19Y5__R2_CONB_0;
  wire tie_lo_T19Y60__R2_CONB_0;
  wire tie_lo_T19Y61__R2_CONB_0;
  wire tie_lo_T19Y62__R2_CONB_0;
  wire tie_lo_T19Y63__R2_CONB_0;
  wire tie_lo_T19Y64__R2_CONB_0;
  wire tie_lo_T19Y65__R2_CONB_0;
  wire tie_lo_T19Y66__R2_CONB_0;
  wire tie_lo_T19Y67__R2_CONB_0;
  wire tie_lo_T19Y68__R2_CONB_0;
  wire tie_lo_T19Y69__R2_CONB_0;
  wire tie_lo_T19Y6__R2_CONB_0;
  wire tie_lo_T19Y70__R2_CONB_0;
  wire tie_lo_T19Y71__R2_CONB_0;
  wire tie_lo_T19Y72__R2_CONB_0;
  wire tie_lo_T19Y73__R2_CONB_0;
  wire tie_lo_T19Y74__R2_CONB_0;
  wire tie_lo_T19Y75__R2_CONB_0;
  wire tie_lo_T19Y76__R2_CONB_0;
  wire tie_lo_T19Y77__R2_CONB_0;
  wire tie_lo_T19Y78__R2_CONB_0;
  wire tie_lo_T19Y79__R2_CONB_0;
  wire tie_lo_T19Y7__R2_CONB_0;
  wire tie_lo_T19Y80__R2_CONB_0;
  wire tie_lo_T19Y81__R2_CONB_0;
  wire tie_lo_T19Y82__R2_CONB_0;
  wire tie_lo_T19Y83__R2_CONB_0;
  wire tie_lo_T19Y84__R2_CONB_0;
  wire tie_lo_T19Y85__R2_CONB_0;
  wire tie_lo_T19Y86__R2_CONB_0;
  wire tie_lo_T19Y87__R2_CONB_0;
  wire tie_lo_T19Y88__R2_CONB_0;
  wire tie_lo_T19Y89__R2_CONB_0;
  wire tie_lo_T19Y8__R2_CONB_0;
  wire tie_lo_T19Y9__R2_CONB_0;
  wire tie_lo_T1Y0__R2_CONB_0;
  wire tie_lo_T1Y10__R2_CONB_0;
  wire tie_lo_T1Y11__R2_CONB_0;
  wire tie_lo_T1Y12__R2_CONB_0;
  wire tie_lo_T1Y13__R2_CONB_0;
  wire tie_lo_T1Y14__R2_CONB_0;
  wire tie_lo_T1Y15__R2_CONB_0;
  wire tie_lo_T1Y16__R2_CONB_0;
  wire tie_lo_T1Y17__R2_CONB_0;
  wire tie_lo_T1Y18__R2_CONB_0;
  wire tie_lo_T1Y19__R2_CONB_0;
  wire tie_lo_T1Y1__R2_CONB_0;
  wire tie_lo_T1Y20__R2_CONB_0;
  wire tie_lo_T1Y21__R2_CONB_0;
  wire tie_lo_T1Y22__R2_CONB_0;
  wire tie_lo_T1Y23__R2_CONB_0;
  wire tie_lo_T1Y24__R2_CONB_0;
  wire tie_lo_T1Y25__R2_CONB_0;
  wire tie_lo_T1Y26__R2_CONB_0;
  wire tie_lo_T1Y27__R2_CONB_0;
  wire tie_lo_T1Y28__R2_CONB_0;
  wire tie_lo_T1Y29__R2_CONB_0;
  wire tie_lo_T1Y2__R2_CONB_0;
  wire tie_lo_T1Y30__R2_CONB_0;
  wire tie_lo_T1Y31__R2_CONB_0;
  wire tie_lo_T1Y32__R2_CONB_0;
  wire tie_lo_T1Y33__R2_CONB_0;
  wire tie_lo_T1Y34__R2_CONB_0;
  wire tie_lo_T1Y35__R2_CONB_0;
  wire tie_lo_T1Y36__R2_CONB_0;
  wire tie_lo_T1Y37__R2_CONB_0;
  wire tie_lo_T1Y38__R2_CONB_0;
  wire tie_lo_T1Y39__R2_CONB_0;
  wire tie_lo_T1Y3__R2_CONB_0;
  wire tie_lo_T1Y40__R2_CONB_0;
  wire tie_lo_T1Y41__R2_CONB_0;
  wire tie_lo_T1Y42__R2_CONB_0;
  wire tie_lo_T1Y43__R2_CONB_0;
  wire tie_lo_T1Y44__R2_CONB_0;
  wire tie_lo_T1Y45__R2_CONB_0;
  wire tie_lo_T1Y46__R2_CONB_0;
  wire tie_lo_T1Y47__R2_CONB_0;
  wire tie_lo_T1Y48__R2_CONB_0;
  wire tie_lo_T1Y49__R2_CONB_0;
  wire tie_lo_T1Y4__R2_CONB_0;
  wire tie_lo_T1Y50__R2_CONB_0;
  wire tie_lo_T1Y51__R2_CONB_0;
  wire tie_lo_T1Y52__R2_CONB_0;
  wire tie_lo_T1Y53__R2_CONB_0;
  wire tie_lo_T1Y54__R2_CONB_0;
  wire tie_lo_T1Y55__R2_CONB_0;
  wire tie_lo_T1Y56__R2_CONB_0;
  wire tie_lo_T1Y57__R2_CONB_0;
  wire tie_lo_T1Y58__R2_CONB_0;
  wire tie_lo_T1Y59__R2_CONB_0;
  wire tie_lo_T1Y5__R2_CONB_0;
  wire tie_lo_T1Y60__R2_CONB_0;
  wire tie_lo_T1Y61__R2_CONB_0;
  wire tie_lo_T1Y62__R2_CONB_0;
  wire tie_lo_T1Y63__R2_CONB_0;
  wire tie_lo_T1Y64__R2_CONB_0;
  wire tie_lo_T1Y65__R2_CONB_0;
  wire tie_lo_T1Y66__R2_CONB_0;
  wire tie_lo_T1Y67__R2_CONB_0;
  wire tie_lo_T1Y68__R2_CONB_0;
  wire tie_lo_T1Y69__R2_CONB_0;
  wire tie_lo_T1Y6__R2_CONB_0;
  wire tie_lo_T1Y70__R2_CONB_0;
  wire tie_lo_T1Y71__R2_CONB_0;
  wire tie_lo_T1Y72__R2_CONB_0;
  wire tie_lo_T1Y73__R2_CONB_0;
  wire tie_lo_T1Y74__R2_CONB_0;
  wire tie_lo_T1Y75__R2_CONB_0;
  wire tie_lo_T1Y76__R2_CONB_0;
  wire tie_lo_T1Y77__R2_CONB_0;
  wire tie_lo_T1Y78__R2_CONB_0;
  wire tie_lo_T1Y79__R2_CONB_0;
  wire tie_lo_T1Y7__R2_CONB_0;
  wire tie_lo_T1Y80__R2_CONB_0;
  wire tie_lo_T1Y81__R2_CONB_0;
  wire tie_lo_T1Y82__R2_CONB_0;
  wire tie_lo_T1Y83__R2_CONB_0;
  wire tie_lo_T1Y84__R2_CONB_0;
  wire tie_lo_T1Y85__R2_CONB_0;
  wire tie_lo_T1Y86__R2_CONB_0;
  wire tie_lo_T1Y87__R2_CONB_0;
  wire tie_lo_T1Y88__R2_CONB_0;
  wire tie_lo_T1Y89__R2_CONB_0;
  wire tie_lo_T1Y8__R2_CONB_0;
  wire tie_lo_T1Y9__R2_CONB_0;
  wire tie_lo_T20Y0__R2_CONB_0;
  wire tie_lo_T20Y10__R2_CONB_0;
  wire tie_lo_T20Y11__R2_CONB_0;
  wire tie_lo_T20Y12__R2_CONB_0;
  wire tie_lo_T20Y13__R2_CONB_0;
  wire tie_lo_T20Y14__R2_CONB_0;
  wire tie_lo_T20Y15__R2_CONB_0;
  wire tie_lo_T20Y16__R2_CONB_0;
  wire tie_lo_T20Y17__R2_CONB_0;
  wire tie_lo_T20Y18__R2_CONB_0;
  wire tie_lo_T20Y19__R2_CONB_0;
  wire tie_lo_T20Y1__R2_CONB_0;
  wire tie_lo_T20Y20__R2_CONB_0;
  wire tie_lo_T20Y21__R2_CONB_0;
  wire tie_lo_T20Y22__R2_CONB_0;
  wire tie_lo_T20Y23__R2_CONB_0;
  wire tie_lo_T20Y24__R2_CONB_0;
  wire tie_lo_T20Y25__R2_CONB_0;
  wire tie_lo_T20Y26__R2_CONB_0;
  wire tie_lo_T20Y27__R2_CONB_0;
  wire tie_lo_T20Y28__R2_CONB_0;
  wire tie_lo_T20Y29__R2_CONB_0;
  wire tie_lo_T20Y2__R2_CONB_0;
  wire tie_lo_T20Y30__R2_CONB_0;
  wire tie_lo_T20Y31__R2_CONB_0;
  wire tie_lo_T20Y32__R2_CONB_0;
  wire tie_lo_T20Y33__R2_CONB_0;
  wire tie_lo_T20Y34__R2_CONB_0;
  wire tie_lo_T20Y35__R2_CONB_0;
  wire tie_lo_T20Y36__R2_CONB_0;
  wire tie_lo_T20Y37__R2_CONB_0;
  wire tie_lo_T20Y38__R2_CONB_0;
  wire tie_lo_T20Y39__R2_CONB_0;
  wire tie_lo_T20Y3__R2_CONB_0;
  wire tie_lo_T20Y40__R2_CONB_0;
  wire tie_lo_T20Y41__R2_CONB_0;
  wire tie_lo_T20Y42__R2_CONB_0;
  wire tie_lo_T20Y43__R2_CONB_0;
  wire tie_lo_T20Y44__R2_CONB_0;
  wire tie_lo_T20Y45__R2_CONB_0;
  wire tie_lo_T20Y46__R2_CONB_0;
  wire tie_lo_T20Y47__R2_CONB_0;
  wire tie_lo_T20Y48__R2_CONB_0;
  wire tie_lo_T20Y49__R2_CONB_0;
  wire tie_lo_T20Y4__R2_CONB_0;
  wire tie_lo_T20Y50__R2_CONB_0;
  wire tie_lo_T20Y51__R2_CONB_0;
  wire tie_lo_T20Y52__R2_CONB_0;
  wire tie_lo_T20Y53__R2_CONB_0;
  wire tie_lo_T20Y54__R2_CONB_0;
  wire tie_lo_T20Y55__R2_CONB_0;
  wire tie_lo_T20Y56__R2_CONB_0;
  wire tie_lo_T20Y57__R2_CONB_0;
  wire tie_lo_T20Y58__R2_CONB_0;
  wire tie_lo_T20Y59__R2_CONB_0;
  wire tie_lo_T20Y5__R2_CONB_0;
  wire tie_lo_T20Y60__R2_CONB_0;
  wire tie_lo_T20Y61__R2_CONB_0;
  wire tie_lo_T20Y62__R2_CONB_0;
  wire tie_lo_T20Y63__R2_CONB_0;
  wire tie_lo_T20Y64__R2_CONB_0;
  wire tie_lo_T20Y65__R2_CONB_0;
  wire tie_lo_T20Y66__R2_CONB_0;
  wire tie_lo_T20Y67__R2_CONB_0;
  wire tie_lo_T20Y68__R2_CONB_0;
  wire tie_lo_T20Y69__R2_CONB_0;
  wire tie_lo_T20Y6__R2_CONB_0;
  wire tie_lo_T20Y70__R2_CONB_0;
  wire tie_lo_T20Y71__R2_CONB_0;
  wire tie_lo_T20Y72__R2_CONB_0;
  wire tie_lo_T20Y73__R2_CONB_0;
  wire tie_lo_T20Y74__R2_CONB_0;
  wire tie_lo_T20Y75__R2_CONB_0;
  wire tie_lo_T20Y76__R2_CONB_0;
  wire tie_lo_T20Y77__R2_CONB_0;
  wire tie_lo_T20Y78__R2_CONB_0;
  wire tie_lo_T20Y79__R2_CONB_0;
  wire tie_lo_T20Y7__R2_CONB_0;
  wire tie_lo_T20Y80__R2_CONB_0;
  wire tie_lo_T20Y81__R2_CONB_0;
  wire tie_lo_T20Y82__R2_CONB_0;
  wire tie_lo_T20Y83__R2_CONB_0;
  wire tie_lo_T20Y84__R2_CONB_0;
  wire tie_lo_T20Y85__R2_CONB_0;
  wire tie_lo_T20Y86__R2_CONB_0;
  wire tie_lo_T20Y87__R2_CONB_0;
  wire tie_lo_T20Y88__R2_CONB_0;
  wire tie_lo_T20Y89__R2_CONB_0;
  wire tie_lo_T20Y8__R2_CONB_0;
  wire tie_lo_T20Y9__R2_CONB_0;
  wire tie_lo_T21Y0__R2_CONB_0;
  wire tie_lo_T21Y10__R2_CONB_0;
  wire tie_lo_T21Y11__R2_CONB_0;
  wire tie_lo_T21Y12__R2_CONB_0;
  wire tie_lo_T21Y13__R2_CONB_0;
  wire tie_lo_T21Y14__R2_CONB_0;
  wire tie_lo_T21Y15__R2_CONB_0;
  wire tie_lo_T21Y16__R2_CONB_0;
  wire tie_lo_T21Y17__R2_CONB_0;
  wire tie_lo_T21Y18__R2_CONB_0;
  wire tie_lo_T21Y19__R2_CONB_0;
  wire tie_lo_T21Y1__R2_CONB_0;
  wire tie_lo_T21Y20__R2_CONB_0;
  wire tie_lo_T21Y21__R2_CONB_0;
  wire tie_lo_T21Y22__R2_CONB_0;
  wire tie_lo_T21Y23__R2_CONB_0;
  wire tie_lo_T21Y24__R2_CONB_0;
  wire tie_lo_T21Y25__R2_CONB_0;
  wire tie_lo_T21Y26__R2_CONB_0;
  wire tie_lo_T21Y27__R2_CONB_0;
  wire tie_lo_T21Y28__R2_CONB_0;
  wire tie_lo_T21Y29__R2_CONB_0;
  wire tie_lo_T21Y2__R2_CONB_0;
  wire tie_lo_T21Y30__R2_CONB_0;
  wire tie_lo_T21Y31__R2_CONB_0;
  wire tie_lo_T21Y32__R2_CONB_0;
  wire tie_lo_T21Y33__R2_CONB_0;
  wire tie_lo_T21Y34__R2_CONB_0;
  wire tie_lo_T21Y35__R2_CONB_0;
  wire tie_lo_T21Y36__R2_CONB_0;
  wire tie_lo_T21Y37__R2_CONB_0;
  wire tie_lo_T21Y38__R2_CONB_0;
  wire tie_lo_T21Y39__R2_CONB_0;
  wire tie_lo_T21Y3__R2_CONB_0;
  wire tie_lo_T21Y40__R2_CONB_0;
  wire tie_lo_T21Y41__R2_CONB_0;
  wire tie_lo_T21Y42__R2_CONB_0;
  wire tie_lo_T21Y43__R2_CONB_0;
  wire tie_lo_T21Y44__R2_CONB_0;
  wire tie_lo_T21Y45__R2_CONB_0;
  wire tie_lo_T21Y46__R2_CONB_0;
  wire tie_lo_T21Y47__R2_CONB_0;
  wire tie_lo_T21Y48__R2_CONB_0;
  wire tie_lo_T21Y49__R2_CONB_0;
  wire tie_lo_T21Y4__R2_CONB_0;
  wire tie_lo_T21Y50__R2_CONB_0;
  wire tie_lo_T21Y51__R2_CONB_0;
  wire tie_lo_T21Y52__R2_CONB_0;
  wire tie_lo_T21Y53__R2_CONB_0;
  wire tie_lo_T21Y54__R2_CONB_0;
  wire tie_lo_T21Y55__R2_CONB_0;
  wire tie_lo_T21Y56__R2_CONB_0;
  wire tie_lo_T21Y57__R2_CONB_0;
  wire tie_lo_T21Y58__R2_CONB_0;
  wire tie_lo_T21Y59__R2_CONB_0;
  wire tie_lo_T21Y5__R2_CONB_0;
  wire tie_lo_T21Y60__R2_CONB_0;
  wire tie_lo_T21Y61__R2_CONB_0;
  wire tie_lo_T21Y62__R2_CONB_0;
  wire tie_lo_T21Y63__R2_CONB_0;
  wire tie_lo_T21Y64__R2_CONB_0;
  wire tie_lo_T21Y65__R2_CONB_0;
  wire tie_lo_T21Y66__R2_CONB_0;
  wire tie_lo_T21Y67__R2_CONB_0;
  wire tie_lo_T21Y68__R2_CONB_0;
  wire tie_lo_T21Y69__R2_CONB_0;
  wire tie_lo_T21Y6__R2_CONB_0;
  wire tie_lo_T21Y70__R2_CONB_0;
  wire tie_lo_T21Y71__R2_CONB_0;
  wire tie_lo_T21Y72__R2_CONB_0;
  wire tie_lo_T21Y73__R2_CONB_0;
  wire tie_lo_T21Y74__R2_CONB_0;
  wire tie_lo_T21Y75__R2_CONB_0;
  wire tie_lo_T21Y76__R2_CONB_0;
  wire tie_lo_T21Y77__R2_CONB_0;
  wire tie_lo_T21Y78__R2_CONB_0;
  wire tie_lo_T21Y79__R2_CONB_0;
  wire tie_lo_T21Y7__R2_CONB_0;
  wire tie_lo_T21Y80__R2_CONB_0;
  wire tie_lo_T21Y81__R2_CONB_0;
  wire tie_lo_T21Y82__R2_CONB_0;
  wire tie_lo_T21Y83__R2_CONB_0;
  wire tie_lo_T21Y84__R2_CONB_0;
  wire tie_lo_T21Y85__R2_CONB_0;
  wire tie_lo_T21Y86__R2_CONB_0;
  wire tie_lo_T21Y87__R2_CONB_0;
  wire tie_lo_T21Y88__R2_CONB_0;
  wire tie_lo_T21Y89__R2_CONB_0;
  wire tie_lo_T21Y8__R2_CONB_0;
  wire tie_lo_T21Y9__R2_CONB_0;
  wire tie_lo_T22Y0__R2_CONB_0;
  wire tie_lo_T22Y10__R2_CONB_0;
  wire tie_lo_T22Y11__R2_CONB_0;
  wire tie_lo_T22Y12__R2_CONB_0;
  wire tie_lo_T22Y13__R2_CONB_0;
  wire tie_lo_T22Y14__R2_CONB_0;
  wire tie_lo_T22Y15__R2_CONB_0;
  wire tie_lo_T22Y16__R2_CONB_0;
  wire tie_lo_T22Y17__R2_CONB_0;
  wire tie_lo_T22Y18__R2_CONB_0;
  wire tie_lo_T22Y19__R2_CONB_0;
  wire tie_lo_T22Y1__R2_CONB_0;
  wire tie_lo_T22Y20__R2_CONB_0;
  wire tie_lo_T22Y21__R2_CONB_0;
  wire tie_lo_T22Y22__R2_CONB_0;
  wire tie_lo_T22Y23__R2_CONB_0;
  wire tie_lo_T22Y24__R2_CONB_0;
  wire tie_lo_T22Y25__R2_CONB_0;
  wire tie_lo_T22Y26__R2_CONB_0;
  wire tie_lo_T22Y27__R2_CONB_0;
  wire tie_lo_T22Y28__R2_CONB_0;
  wire tie_lo_T22Y29__R2_CONB_0;
  wire tie_lo_T22Y2__R2_CONB_0;
  wire tie_lo_T22Y30__R2_CONB_0;
  wire tie_lo_T22Y31__R2_CONB_0;
  wire tie_lo_T22Y32__R2_CONB_0;
  wire tie_lo_T22Y33__R2_CONB_0;
  wire tie_lo_T22Y34__R2_CONB_0;
  wire tie_lo_T22Y35__R2_CONB_0;
  wire tie_lo_T22Y36__R2_CONB_0;
  wire tie_lo_T22Y37__R2_CONB_0;
  wire tie_lo_T22Y38__R2_CONB_0;
  wire tie_lo_T22Y39__R2_CONB_0;
  wire tie_lo_T22Y3__R2_CONB_0;
  wire tie_lo_T22Y40__R2_CONB_0;
  wire tie_lo_T22Y41__R2_CONB_0;
  wire tie_lo_T22Y42__R2_CONB_0;
  wire tie_lo_T22Y43__R2_CONB_0;
  wire tie_lo_T22Y44__R2_CONB_0;
  wire tie_lo_T22Y45__R2_CONB_0;
  wire tie_lo_T22Y46__R2_CONB_0;
  wire tie_lo_T22Y47__R2_CONB_0;
  wire tie_lo_T22Y48__R2_CONB_0;
  wire tie_lo_T22Y49__R2_CONB_0;
  wire tie_lo_T22Y4__R2_CONB_0;
  wire tie_lo_T22Y50__R2_CONB_0;
  wire tie_lo_T22Y51__R2_CONB_0;
  wire tie_lo_T22Y52__R2_CONB_0;
  wire tie_lo_T22Y53__R2_CONB_0;
  wire tie_lo_T22Y54__R2_CONB_0;
  wire tie_lo_T22Y55__R2_CONB_0;
  wire tie_lo_T22Y56__R2_CONB_0;
  wire tie_lo_T22Y57__R2_CONB_0;
  wire tie_lo_T22Y58__R2_CONB_0;
  wire tie_lo_T22Y59__R2_CONB_0;
  wire tie_lo_T22Y5__R2_CONB_0;
  wire tie_lo_T22Y60__R2_CONB_0;
  wire tie_lo_T22Y61__R2_CONB_0;
  wire tie_lo_T22Y62__R2_CONB_0;
  wire tie_lo_T22Y63__R2_CONB_0;
  wire tie_lo_T22Y64__R2_CONB_0;
  wire tie_lo_T22Y65__R2_CONB_0;
  wire tie_lo_T22Y66__R2_CONB_0;
  wire tie_lo_T22Y67__R2_CONB_0;
  wire tie_lo_T22Y68__R2_CONB_0;
  wire tie_lo_T22Y69__R2_CONB_0;
  wire tie_lo_T22Y6__R2_CONB_0;
  wire tie_lo_T22Y70__R2_CONB_0;
  wire tie_lo_T22Y71__R2_CONB_0;
  wire tie_lo_T22Y72__R2_CONB_0;
  wire tie_lo_T22Y73__R2_CONB_0;
  wire tie_lo_T22Y74__R2_CONB_0;
  wire tie_lo_T22Y75__R2_CONB_0;
  wire tie_lo_T22Y76__R2_CONB_0;
  wire tie_lo_T22Y77__R2_CONB_0;
  wire tie_lo_T22Y78__R2_CONB_0;
  wire tie_lo_T22Y79__R2_CONB_0;
  wire tie_lo_T22Y7__R2_CONB_0;
  wire tie_lo_T22Y80__R2_CONB_0;
  wire tie_lo_T22Y81__R2_CONB_0;
  wire tie_lo_T22Y82__R2_CONB_0;
  wire tie_lo_T22Y83__R2_CONB_0;
  wire tie_lo_T22Y84__R2_CONB_0;
  wire tie_lo_T22Y85__R2_CONB_0;
  wire tie_lo_T22Y86__R2_CONB_0;
  wire tie_lo_T22Y87__R2_CONB_0;
  wire tie_lo_T22Y88__R2_CONB_0;
  wire tie_lo_T22Y89__R2_CONB_0;
  wire tie_lo_T22Y8__R2_CONB_0;
  wire tie_lo_T22Y9__R2_CONB_0;
  wire tie_lo_T23Y0__R2_CONB_0;
  wire tie_lo_T23Y10__R2_CONB_0;
  wire tie_lo_T23Y11__R2_CONB_0;
  wire tie_lo_T23Y12__R2_CONB_0;
  wire tie_lo_T23Y13__R2_CONB_0;
  wire tie_lo_T23Y14__R2_CONB_0;
  wire tie_lo_T23Y15__R2_CONB_0;
  wire tie_lo_T23Y16__R2_CONB_0;
  wire tie_lo_T23Y17__R2_CONB_0;
  wire tie_lo_T23Y18__R2_CONB_0;
  wire tie_lo_T23Y19__R2_CONB_0;
  wire tie_lo_T23Y1__R2_CONB_0;
  wire tie_lo_T23Y20__R2_CONB_0;
  wire tie_lo_T23Y21__R2_CONB_0;
  wire tie_lo_T23Y22__R2_CONB_0;
  wire tie_lo_T23Y23__R2_CONB_0;
  wire tie_lo_T23Y24__R2_CONB_0;
  wire tie_lo_T23Y25__R2_CONB_0;
  wire tie_lo_T23Y26__R2_CONB_0;
  wire tie_lo_T23Y27__R2_CONB_0;
  wire tie_lo_T23Y28__R2_CONB_0;
  wire tie_lo_T23Y29__R2_CONB_0;
  wire tie_lo_T23Y2__R2_CONB_0;
  wire tie_lo_T23Y30__R2_CONB_0;
  wire tie_lo_T23Y31__R2_CONB_0;
  wire tie_lo_T23Y32__R2_CONB_0;
  wire tie_lo_T23Y33__R2_CONB_0;
  wire tie_lo_T23Y34__R2_CONB_0;
  wire tie_lo_T23Y35__R2_CONB_0;
  wire tie_lo_T23Y36__R2_CONB_0;
  wire tie_lo_T23Y37__R2_CONB_0;
  wire tie_lo_T23Y38__R2_CONB_0;
  wire tie_lo_T23Y39__R2_CONB_0;
  wire tie_lo_T23Y3__R2_CONB_0;
  wire tie_lo_T23Y40__R2_CONB_0;
  wire tie_lo_T23Y41__R2_CONB_0;
  wire tie_lo_T23Y42__R2_CONB_0;
  wire tie_lo_T23Y43__R2_CONB_0;
  wire tie_lo_T23Y44__R2_CONB_0;
  wire tie_lo_T23Y45__R2_CONB_0;
  wire tie_lo_T23Y46__R2_CONB_0;
  wire tie_lo_T23Y47__R2_CONB_0;
  wire tie_lo_T23Y48__R2_CONB_0;
  wire tie_lo_T23Y49__R2_CONB_0;
  wire tie_lo_T23Y4__R2_CONB_0;
  wire tie_lo_T23Y50__R2_CONB_0;
  wire tie_lo_T23Y51__R2_CONB_0;
  wire tie_lo_T23Y52__R2_CONB_0;
  wire tie_lo_T23Y53__R2_CONB_0;
  wire tie_lo_T23Y54__R2_CONB_0;
  wire tie_lo_T23Y55__R2_CONB_0;
  wire tie_lo_T23Y56__R2_CONB_0;
  wire tie_lo_T23Y57__R2_CONB_0;
  wire tie_lo_T23Y58__R2_CONB_0;
  wire tie_lo_T23Y59__R2_CONB_0;
  wire tie_lo_T23Y5__R2_CONB_0;
  wire tie_lo_T23Y60__R2_CONB_0;
  wire tie_lo_T23Y61__R2_CONB_0;
  wire tie_lo_T23Y62__R2_CONB_0;
  wire tie_lo_T23Y63__R2_CONB_0;
  wire tie_lo_T23Y64__R2_CONB_0;
  wire tie_lo_T23Y65__R2_CONB_0;
  wire tie_lo_T23Y66__R2_CONB_0;
  wire tie_lo_T23Y67__R2_CONB_0;
  wire tie_lo_T23Y68__R2_CONB_0;
  wire tie_lo_T23Y69__R2_CONB_0;
  wire tie_lo_T23Y6__R2_CONB_0;
  wire tie_lo_T23Y70__R2_CONB_0;
  wire tie_lo_T23Y71__R2_CONB_0;
  wire tie_lo_T23Y72__R2_CONB_0;
  wire tie_lo_T23Y73__R2_CONB_0;
  wire tie_lo_T23Y74__R2_CONB_0;
  wire tie_lo_T23Y75__R2_CONB_0;
  wire tie_lo_T23Y76__R2_CONB_0;
  wire tie_lo_T23Y77__R2_CONB_0;
  wire tie_lo_T23Y78__R2_CONB_0;
  wire tie_lo_T23Y79__R2_CONB_0;
  wire tie_lo_T23Y7__R2_CONB_0;
  wire tie_lo_T23Y80__R2_CONB_0;
  wire tie_lo_T23Y81__R2_CONB_0;
  wire tie_lo_T23Y82__R2_CONB_0;
  wire tie_lo_T23Y83__R2_CONB_0;
  wire tie_lo_T23Y84__R2_CONB_0;
  wire tie_lo_T23Y85__R2_CONB_0;
  wire tie_lo_T23Y86__R2_CONB_0;
  wire tie_lo_T23Y87__R2_CONB_0;
  wire tie_lo_T23Y88__R2_CONB_0;
  wire tie_lo_T23Y89__R2_CONB_0;
  wire tie_lo_T23Y8__R2_CONB_0;
  wire tie_lo_T23Y9__R2_CONB_0;
  wire tie_lo_T24Y0__R2_CONB_0;
  wire tie_lo_T24Y10__R2_CONB_0;
  wire tie_lo_T24Y11__R2_CONB_0;
  wire tie_lo_T24Y12__R2_CONB_0;
  wire tie_lo_T24Y13__R2_CONB_0;
  wire tie_lo_T24Y14__R2_CONB_0;
  wire tie_lo_T24Y15__R2_CONB_0;
  wire tie_lo_T24Y16__R2_CONB_0;
  wire tie_lo_T24Y17__R2_CONB_0;
  wire tie_lo_T24Y18__R2_CONB_0;
  wire tie_lo_T24Y19__R2_CONB_0;
  wire tie_lo_T24Y1__R2_CONB_0;
  wire tie_lo_T24Y20__R2_CONB_0;
  wire tie_lo_T24Y21__R2_CONB_0;
  wire tie_lo_T24Y22__R2_CONB_0;
  wire tie_lo_T24Y23__R2_CONB_0;
  wire tie_lo_T24Y24__R2_CONB_0;
  wire tie_lo_T24Y25__R2_CONB_0;
  wire tie_lo_T24Y26__R2_CONB_0;
  wire tie_lo_T24Y27__R2_CONB_0;
  wire tie_lo_T24Y28__R2_CONB_0;
  wire tie_lo_T24Y29__R2_CONB_0;
  wire tie_lo_T24Y2__R2_CONB_0;
  wire tie_lo_T24Y30__R2_CONB_0;
  wire tie_lo_T24Y31__R2_CONB_0;
  wire tie_lo_T24Y32__R2_CONB_0;
  wire tie_lo_T24Y33__R2_CONB_0;
  wire tie_lo_T24Y34__R2_CONB_0;
  wire tie_lo_T24Y35__R2_CONB_0;
  wire tie_lo_T24Y36__R2_CONB_0;
  wire tie_lo_T24Y37__R2_CONB_0;
  wire tie_lo_T24Y38__R2_CONB_0;
  wire tie_lo_T24Y39__R2_CONB_0;
  wire tie_lo_T24Y3__R2_CONB_0;
  wire tie_lo_T24Y40__R2_CONB_0;
  wire tie_lo_T24Y41__R2_CONB_0;
  wire tie_lo_T24Y42__R2_CONB_0;
  wire tie_lo_T24Y43__R2_CONB_0;
  wire tie_lo_T24Y44__R2_CONB_0;
  wire tie_lo_T24Y45__R2_CONB_0;
  wire tie_lo_T24Y46__R2_CONB_0;
  wire tie_lo_T24Y47__R2_CONB_0;
  wire tie_lo_T24Y48__R2_CONB_0;
  wire tie_lo_T24Y49__R2_CONB_0;
  wire tie_lo_T24Y4__R2_CONB_0;
  wire tie_lo_T24Y50__R2_CONB_0;
  wire tie_lo_T24Y51__R2_CONB_0;
  wire tie_lo_T24Y52__R2_CONB_0;
  wire tie_lo_T24Y53__R2_CONB_0;
  wire tie_lo_T24Y54__R2_CONB_0;
  wire tie_lo_T24Y55__R2_CONB_0;
  wire tie_lo_T24Y56__R2_CONB_0;
  wire tie_lo_T24Y57__R2_CONB_0;
  wire tie_lo_T24Y58__R2_CONB_0;
  wire tie_lo_T24Y59__R2_CONB_0;
  wire tie_lo_T24Y5__R2_CONB_0;
  wire tie_lo_T24Y60__R2_CONB_0;
  wire tie_lo_T24Y61__R2_CONB_0;
  wire tie_lo_T24Y62__R2_CONB_0;
  wire tie_lo_T24Y63__R2_CONB_0;
  wire tie_lo_T24Y64__R2_CONB_0;
  wire tie_lo_T24Y65__R2_CONB_0;
  wire tie_lo_T24Y66__R2_CONB_0;
  wire tie_lo_T24Y67__R2_CONB_0;
  wire tie_lo_T24Y68__R2_CONB_0;
  wire tie_lo_T24Y69__R2_CONB_0;
  wire tie_lo_T24Y6__R2_CONB_0;
  wire tie_lo_T24Y70__R2_CONB_0;
  wire tie_lo_T24Y71__R2_CONB_0;
  wire tie_lo_T24Y72__R2_CONB_0;
  wire tie_lo_T24Y73__R2_CONB_0;
  wire tie_lo_T24Y74__R2_CONB_0;
  wire tie_lo_T24Y75__R2_CONB_0;
  wire tie_lo_T24Y76__R2_CONB_0;
  wire tie_lo_T24Y77__R2_CONB_0;
  wire tie_lo_T24Y78__R2_CONB_0;
  wire tie_lo_T24Y79__R2_CONB_0;
  wire tie_lo_T24Y7__R2_CONB_0;
  wire tie_lo_T24Y80__R2_CONB_0;
  wire tie_lo_T24Y81__R2_CONB_0;
  wire tie_lo_T24Y82__R2_CONB_0;
  wire tie_lo_T24Y83__R2_CONB_0;
  wire tie_lo_T24Y84__R2_CONB_0;
  wire tie_lo_T24Y85__R2_CONB_0;
  wire tie_lo_T24Y86__R2_CONB_0;
  wire tie_lo_T24Y87__R2_CONB_0;
  wire tie_lo_T24Y88__R2_CONB_0;
  wire tie_lo_T24Y89__R2_CONB_0;
  wire tie_lo_T24Y8__R2_CONB_0;
  wire tie_lo_T24Y9__R2_CONB_0;
  wire tie_lo_T25Y0__R2_CONB_0;
  wire tie_lo_T25Y10__R2_CONB_0;
  wire tie_lo_T25Y11__R2_CONB_0;
  wire tie_lo_T25Y12__R2_CONB_0;
  wire tie_lo_T25Y13__R2_CONB_0;
  wire tie_lo_T25Y14__R2_CONB_0;
  wire tie_lo_T25Y15__R2_CONB_0;
  wire tie_lo_T25Y16__R2_CONB_0;
  wire tie_lo_T25Y17__R2_CONB_0;
  wire tie_lo_T25Y18__R2_CONB_0;
  wire tie_lo_T25Y19__R2_CONB_0;
  wire tie_lo_T25Y1__R2_CONB_0;
  wire tie_lo_T25Y20__R2_CONB_0;
  wire tie_lo_T25Y21__R2_CONB_0;
  wire tie_lo_T25Y22__R2_CONB_0;
  wire tie_lo_T25Y23__R2_CONB_0;
  wire tie_lo_T25Y24__R2_CONB_0;
  wire tie_lo_T25Y25__R2_CONB_0;
  wire tie_lo_T25Y26__R2_CONB_0;
  wire tie_lo_T25Y27__R2_CONB_0;
  wire tie_lo_T25Y28__R2_CONB_0;
  wire tie_lo_T25Y29__R2_CONB_0;
  wire tie_lo_T25Y2__R2_CONB_0;
  wire tie_lo_T25Y30__R2_CONB_0;
  wire tie_lo_T25Y31__R2_CONB_0;
  wire tie_lo_T25Y32__R2_CONB_0;
  wire tie_lo_T25Y33__R2_CONB_0;
  wire tie_lo_T25Y34__R2_CONB_0;
  wire tie_lo_T25Y35__R2_CONB_0;
  wire tie_lo_T25Y36__R2_CONB_0;
  wire tie_lo_T25Y37__R2_CONB_0;
  wire tie_lo_T25Y38__R2_CONB_0;
  wire tie_lo_T25Y39__R2_CONB_0;
  wire tie_lo_T25Y3__R2_CONB_0;
  wire tie_lo_T25Y40__R2_CONB_0;
  wire tie_lo_T25Y41__R2_CONB_0;
  wire tie_lo_T25Y42__R2_CONB_0;
  wire tie_lo_T25Y43__R2_CONB_0;
  wire tie_lo_T25Y44__R2_CONB_0;
  wire tie_lo_T25Y45__R2_CONB_0;
  wire tie_lo_T25Y46__R2_CONB_0;
  wire tie_lo_T25Y47__R2_CONB_0;
  wire tie_lo_T25Y48__R2_CONB_0;
  wire tie_lo_T25Y49__R2_CONB_0;
  wire tie_lo_T25Y4__R2_CONB_0;
  wire tie_lo_T25Y50__R2_CONB_0;
  wire tie_lo_T25Y51__R2_CONB_0;
  wire tie_lo_T25Y52__R2_CONB_0;
  wire tie_lo_T25Y53__R2_CONB_0;
  wire tie_lo_T25Y54__R2_CONB_0;
  wire tie_lo_T25Y55__R2_CONB_0;
  wire tie_lo_T25Y56__R2_CONB_0;
  wire tie_lo_T25Y57__R2_CONB_0;
  wire tie_lo_T25Y58__R2_CONB_0;
  wire tie_lo_T25Y59__R2_CONB_0;
  wire tie_lo_T25Y5__R2_CONB_0;
  wire tie_lo_T25Y60__R2_CONB_0;
  wire tie_lo_T25Y61__R2_CONB_0;
  wire tie_lo_T25Y62__R2_CONB_0;
  wire tie_lo_T25Y63__R2_CONB_0;
  wire tie_lo_T25Y64__R2_CONB_0;
  wire tie_lo_T25Y65__R2_CONB_0;
  wire tie_lo_T25Y66__R2_CONB_0;
  wire tie_lo_T25Y67__R2_CONB_0;
  wire tie_lo_T25Y68__R2_CONB_0;
  wire tie_lo_T25Y69__R2_CONB_0;
  wire tie_lo_T25Y6__R2_CONB_0;
  wire tie_lo_T25Y70__R2_CONB_0;
  wire tie_lo_T25Y71__R2_CONB_0;
  wire tie_lo_T25Y72__R2_CONB_0;
  wire tie_lo_T25Y73__R2_CONB_0;
  wire tie_lo_T25Y74__R2_CONB_0;
  wire tie_lo_T25Y75__R2_CONB_0;
  wire tie_lo_T25Y76__R2_CONB_0;
  wire tie_lo_T25Y77__R2_CONB_0;
  wire tie_lo_T25Y78__R2_CONB_0;
  wire tie_lo_T25Y79__R2_CONB_0;
  wire tie_lo_T25Y7__R2_CONB_0;
  wire tie_lo_T25Y80__R2_CONB_0;
  wire tie_lo_T25Y81__R2_CONB_0;
  wire tie_lo_T25Y82__R2_CONB_0;
  wire tie_lo_T25Y83__R2_CONB_0;
  wire tie_lo_T25Y84__R2_CONB_0;
  wire tie_lo_T25Y85__R2_CONB_0;
  wire tie_lo_T25Y86__R2_CONB_0;
  wire tie_lo_T25Y87__R2_CONB_0;
  wire tie_lo_T25Y88__R2_CONB_0;
  wire tie_lo_T25Y89__R2_CONB_0;
  wire tie_lo_T25Y8__R2_CONB_0;
  wire tie_lo_T25Y9__R2_CONB_0;
  wire tie_lo_T26Y0__R2_CONB_0;
  wire tie_lo_T26Y10__R2_CONB_0;
  wire tie_lo_T26Y11__R2_CONB_0;
  wire tie_lo_T26Y12__R2_CONB_0;
  wire tie_lo_T26Y13__R2_CONB_0;
  wire tie_lo_T26Y14__R2_CONB_0;
  wire tie_lo_T26Y15__R2_CONB_0;
  wire tie_lo_T26Y16__R2_CONB_0;
  wire tie_lo_T26Y17__R2_CONB_0;
  wire tie_lo_T26Y18__R2_CONB_0;
  wire tie_lo_T26Y19__R2_CONB_0;
  wire tie_lo_T26Y1__R2_CONB_0;
  wire tie_lo_T26Y20__R2_CONB_0;
  wire tie_lo_T26Y21__R2_CONB_0;
  wire tie_lo_T26Y22__R2_CONB_0;
  wire tie_lo_T26Y23__R2_CONB_0;
  wire tie_lo_T26Y24__R2_CONB_0;
  wire tie_lo_T26Y25__R2_CONB_0;
  wire tie_lo_T26Y26__R2_CONB_0;
  wire tie_lo_T26Y27__R2_CONB_0;
  wire tie_lo_T26Y28__R2_CONB_0;
  wire tie_lo_T26Y29__R2_CONB_0;
  wire tie_lo_T26Y2__R2_CONB_0;
  wire tie_lo_T26Y30__R2_CONB_0;
  wire tie_lo_T26Y31__R2_CONB_0;
  wire tie_lo_T26Y32__R2_CONB_0;
  wire tie_lo_T26Y33__R2_CONB_0;
  wire tie_lo_T26Y34__R2_CONB_0;
  wire tie_lo_T26Y35__R2_CONB_0;
  wire tie_lo_T26Y36__R2_CONB_0;
  wire tie_lo_T26Y37__R2_CONB_0;
  wire tie_lo_T26Y38__R2_CONB_0;
  wire tie_lo_T26Y39__R2_CONB_0;
  wire tie_lo_T26Y3__R2_CONB_0;
  wire tie_lo_T26Y40__R2_CONB_0;
  wire tie_lo_T26Y41__R2_CONB_0;
  wire tie_lo_T26Y42__R2_CONB_0;
  wire tie_lo_T26Y43__R2_CONB_0;
  wire tie_lo_T26Y44__R2_CONB_0;
  wire tie_lo_T26Y45__R2_CONB_0;
  wire tie_lo_T26Y46__R2_CONB_0;
  wire tie_lo_T26Y47__R2_CONB_0;
  wire tie_lo_T26Y48__R2_CONB_0;
  wire tie_lo_T26Y49__R2_CONB_0;
  wire tie_lo_T26Y4__R2_CONB_0;
  wire tie_lo_T26Y50__R2_CONB_0;
  wire tie_lo_T26Y51__R2_CONB_0;
  wire tie_lo_T26Y52__R2_CONB_0;
  wire tie_lo_T26Y53__R2_CONB_0;
  wire tie_lo_T26Y54__R2_CONB_0;
  wire tie_lo_T26Y55__R2_CONB_0;
  wire tie_lo_T26Y56__R2_CONB_0;
  wire tie_lo_T26Y57__R2_CONB_0;
  wire tie_lo_T26Y58__R2_CONB_0;
  wire tie_lo_T26Y59__R2_CONB_0;
  wire tie_lo_T26Y5__R2_CONB_0;
  wire tie_lo_T26Y60__R2_CONB_0;
  wire tie_lo_T26Y61__R2_CONB_0;
  wire tie_lo_T26Y62__R2_CONB_0;
  wire tie_lo_T26Y63__R2_CONB_0;
  wire tie_lo_T26Y64__R2_CONB_0;
  wire tie_lo_T26Y65__R2_CONB_0;
  wire tie_lo_T26Y66__R2_CONB_0;
  wire tie_lo_T26Y67__R2_CONB_0;
  wire tie_lo_T26Y68__R2_CONB_0;
  wire tie_lo_T26Y69__R2_CONB_0;
  wire tie_lo_T26Y6__R2_CONB_0;
  wire tie_lo_T26Y70__R2_CONB_0;
  wire tie_lo_T26Y71__R2_CONB_0;
  wire tie_lo_T26Y72__R2_CONB_0;
  wire tie_lo_T26Y73__R2_CONB_0;
  wire tie_lo_T26Y74__R2_CONB_0;
  wire tie_lo_T26Y75__R2_CONB_0;
  wire tie_lo_T26Y76__R2_CONB_0;
  wire tie_lo_T26Y77__R2_CONB_0;
  wire tie_lo_T26Y78__R2_CONB_0;
  wire tie_lo_T26Y79__R2_CONB_0;
  wire tie_lo_T26Y7__R2_CONB_0;
  wire tie_lo_T26Y80__R2_CONB_0;
  wire tie_lo_T26Y81__R2_CONB_0;
  wire tie_lo_T26Y82__R2_CONB_0;
  wire tie_lo_T26Y83__R2_CONB_0;
  wire tie_lo_T26Y84__R2_CONB_0;
  wire tie_lo_T26Y85__R2_CONB_0;
  wire tie_lo_T26Y86__R2_CONB_0;
  wire tie_lo_T26Y87__R2_CONB_0;
  wire tie_lo_T26Y88__R2_CONB_0;
  wire tie_lo_T26Y89__R2_CONB_0;
  wire tie_lo_T26Y8__R2_CONB_0;
  wire tie_lo_T26Y9__R2_CONB_0;
  wire tie_lo_T27Y0__R2_CONB_0;
  wire tie_lo_T27Y10__R2_CONB_0;
  wire tie_lo_T27Y11__R2_CONB_0;
  wire tie_lo_T27Y12__R2_CONB_0;
  wire tie_lo_T27Y13__R2_CONB_0;
  wire tie_lo_T27Y14__R2_CONB_0;
  wire tie_lo_T27Y15__R2_CONB_0;
  wire tie_lo_T27Y16__R2_CONB_0;
  wire tie_lo_T27Y17__R2_CONB_0;
  wire tie_lo_T27Y18__R2_CONB_0;
  wire tie_lo_T27Y19__R2_CONB_0;
  wire tie_lo_T27Y1__R2_CONB_0;
  wire tie_lo_T27Y20__R2_CONB_0;
  wire tie_lo_T27Y21__R2_CONB_0;
  wire tie_lo_T27Y22__R2_CONB_0;
  wire tie_lo_T27Y23__R2_CONB_0;
  wire tie_lo_T27Y24__R2_CONB_0;
  wire tie_lo_T27Y25__R2_CONB_0;
  wire tie_lo_T27Y26__R2_CONB_0;
  wire tie_lo_T27Y27__R2_CONB_0;
  wire tie_lo_T27Y28__R2_CONB_0;
  wire tie_lo_T27Y29__R2_CONB_0;
  wire tie_lo_T27Y2__R2_CONB_0;
  wire tie_lo_T27Y30__R2_CONB_0;
  wire tie_lo_T27Y31__R2_CONB_0;
  wire tie_lo_T27Y32__R2_CONB_0;
  wire tie_lo_T27Y33__R2_CONB_0;
  wire tie_lo_T27Y34__R2_CONB_0;
  wire tie_lo_T27Y35__R2_CONB_0;
  wire tie_lo_T27Y36__R2_CONB_0;
  wire tie_lo_T27Y37__R2_CONB_0;
  wire tie_lo_T27Y38__R2_CONB_0;
  wire tie_lo_T27Y39__R2_CONB_0;
  wire tie_lo_T27Y3__R2_CONB_0;
  wire tie_lo_T27Y40__R2_CONB_0;
  wire tie_lo_T27Y41__R2_CONB_0;
  wire tie_lo_T27Y42__R2_CONB_0;
  wire tie_lo_T27Y43__R2_CONB_0;
  wire tie_lo_T27Y44__R2_CONB_0;
  wire tie_lo_T27Y45__R2_CONB_0;
  wire tie_lo_T27Y46__R2_CONB_0;
  wire tie_lo_T27Y47__R2_CONB_0;
  wire tie_lo_T27Y48__R2_CONB_0;
  wire tie_lo_T27Y49__R2_CONB_0;
  wire tie_lo_T27Y4__R2_CONB_0;
  wire tie_lo_T27Y50__R2_CONB_0;
  wire tie_lo_T27Y51__R2_CONB_0;
  wire tie_lo_T27Y52__R2_CONB_0;
  wire tie_lo_T27Y53__R2_CONB_0;
  wire tie_lo_T27Y54__R2_CONB_0;
  wire tie_lo_T27Y55__R2_CONB_0;
  wire tie_lo_T27Y56__R2_CONB_0;
  wire tie_lo_T27Y57__R2_CONB_0;
  wire tie_lo_T27Y58__R2_CONB_0;
  wire tie_lo_T27Y59__R2_CONB_0;
  wire tie_lo_T27Y5__R2_CONB_0;
  wire tie_lo_T27Y60__R2_CONB_0;
  wire tie_lo_T27Y61__R2_CONB_0;
  wire tie_lo_T27Y62__R2_CONB_0;
  wire tie_lo_T27Y63__R2_CONB_0;
  wire tie_lo_T27Y64__R2_CONB_0;
  wire tie_lo_T27Y65__R2_CONB_0;
  wire tie_lo_T27Y66__R2_CONB_0;
  wire tie_lo_T27Y67__R2_CONB_0;
  wire tie_lo_T27Y68__R2_CONB_0;
  wire tie_lo_T27Y69__R2_CONB_0;
  wire tie_lo_T27Y6__R2_CONB_0;
  wire tie_lo_T27Y70__R2_CONB_0;
  wire tie_lo_T27Y71__R2_CONB_0;
  wire tie_lo_T27Y72__R2_CONB_0;
  wire tie_lo_T27Y73__R2_CONB_0;
  wire tie_lo_T27Y74__R2_CONB_0;
  wire tie_lo_T27Y75__R2_CONB_0;
  wire tie_lo_T27Y76__R2_CONB_0;
  wire tie_lo_T27Y77__R2_CONB_0;
  wire tie_lo_T27Y78__R2_CONB_0;
  wire tie_lo_T27Y79__R2_CONB_0;
  wire tie_lo_T27Y7__R2_CONB_0;
  wire tie_lo_T27Y80__R2_CONB_0;
  wire tie_lo_T27Y81__R2_CONB_0;
  wire tie_lo_T27Y82__R2_CONB_0;
  wire tie_lo_T27Y83__R2_CONB_0;
  wire tie_lo_T27Y84__R2_CONB_0;
  wire tie_lo_T27Y85__R2_CONB_0;
  wire tie_lo_T27Y86__R2_CONB_0;
  wire tie_lo_T27Y87__R2_CONB_0;
  wire tie_lo_T27Y88__R2_CONB_0;
  wire tie_lo_T27Y89__R2_CONB_0;
  wire tie_lo_T27Y8__R2_CONB_0;
  wire tie_lo_T27Y9__R2_CONB_0;
  wire tie_lo_T28Y0__R2_CONB_0;
  wire tie_lo_T28Y10__R2_CONB_0;
  wire tie_lo_T28Y11__R2_CONB_0;
  wire tie_lo_T28Y12__R2_CONB_0;
  wire tie_lo_T28Y13__R2_CONB_0;
  wire tie_lo_T28Y14__R2_CONB_0;
  wire tie_lo_T28Y15__R2_CONB_0;
  wire tie_lo_T28Y16__R2_CONB_0;
  wire tie_lo_T28Y17__R2_CONB_0;
  wire tie_lo_T28Y18__R2_CONB_0;
  wire tie_lo_T28Y19__R2_CONB_0;
  wire tie_lo_T28Y1__R2_CONB_0;
  wire tie_lo_T28Y20__R2_CONB_0;
  wire tie_lo_T28Y21__R2_CONB_0;
  wire tie_lo_T28Y22__R2_CONB_0;
  wire tie_lo_T28Y23__R2_CONB_0;
  wire tie_lo_T28Y24__R2_CONB_0;
  wire tie_lo_T28Y25__R2_CONB_0;
  wire tie_lo_T28Y26__R2_CONB_0;
  wire tie_lo_T28Y27__R2_CONB_0;
  wire tie_lo_T28Y28__R2_CONB_0;
  wire tie_lo_T28Y29__R2_CONB_0;
  wire tie_lo_T28Y2__R2_CONB_0;
  wire tie_lo_T28Y30__R2_CONB_0;
  wire tie_lo_T28Y31__R2_CONB_0;
  wire tie_lo_T28Y32__R2_CONB_0;
  wire tie_lo_T28Y33__R2_CONB_0;
  wire tie_lo_T28Y34__R2_CONB_0;
  wire tie_lo_T28Y35__R2_CONB_0;
  wire tie_lo_T28Y36__R2_CONB_0;
  wire tie_lo_T28Y37__R2_CONB_0;
  wire tie_lo_T28Y38__R2_CONB_0;
  wire tie_lo_T28Y39__R2_CONB_0;
  wire tie_lo_T28Y3__R2_CONB_0;
  wire tie_lo_T28Y40__R2_CONB_0;
  wire tie_lo_T28Y41__R2_CONB_0;
  wire tie_lo_T28Y42__R2_CONB_0;
  wire tie_lo_T28Y43__R2_CONB_0;
  wire tie_lo_T28Y44__R2_CONB_0;
  wire tie_lo_T28Y45__R2_CONB_0;
  wire tie_lo_T28Y46__R2_CONB_0;
  wire tie_lo_T28Y47__R2_CONB_0;
  wire tie_lo_T28Y48__R2_CONB_0;
  wire tie_lo_T28Y49__R2_CONB_0;
  wire tie_lo_T28Y4__R2_CONB_0;
  wire tie_lo_T28Y50__R2_CONB_0;
  wire tie_lo_T28Y51__R2_CONB_0;
  wire tie_lo_T28Y52__R2_CONB_0;
  wire tie_lo_T28Y53__R2_CONB_0;
  wire tie_lo_T28Y54__R2_CONB_0;
  wire tie_lo_T28Y55__R2_CONB_0;
  wire tie_lo_T28Y56__R2_CONB_0;
  wire tie_lo_T28Y57__R2_CONB_0;
  wire tie_lo_T28Y58__R2_CONB_0;
  wire tie_lo_T28Y59__R2_CONB_0;
  wire tie_lo_T28Y5__R2_CONB_0;
  wire tie_lo_T28Y60__R2_CONB_0;
  wire tie_lo_T28Y61__R2_CONB_0;
  wire tie_lo_T28Y62__R2_CONB_0;
  wire tie_lo_T28Y63__R2_CONB_0;
  wire tie_lo_T28Y64__R2_CONB_0;
  wire tie_lo_T28Y65__R2_CONB_0;
  wire tie_lo_T28Y66__R2_CONB_0;
  wire tie_lo_T28Y67__R2_CONB_0;
  wire tie_lo_T28Y68__R2_CONB_0;
  wire tie_lo_T28Y69__R2_CONB_0;
  wire tie_lo_T28Y6__R2_CONB_0;
  wire tie_lo_T28Y70__R2_CONB_0;
  wire tie_lo_T28Y71__R2_CONB_0;
  wire tie_lo_T28Y72__R2_CONB_0;
  wire tie_lo_T28Y73__R2_CONB_0;
  wire tie_lo_T28Y74__R2_CONB_0;
  wire tie_lo_T28Y75__R2_CONB_0;
  wire tie_lo_T28Y76__R2_CONB_0;
  wire tie_lo_T28Y77__R2_CONB_0;
  wire tie_lo_T28Y78__R2_CONB_0;
  wire tie_lo_T28Y79__R2_CONB_0;
  wire tie_lo_T28Y7__R2_CONB_0;
  wire tie_lo_T28Y80__R2_CONB_0;
  wire tie_lo_T28Y81__R2_CONB_0;
  wire tie_lo_T28Y82__R2_CONB_0;
  wire tie_lo_T28Y83__R2_CONB_0;
  wire tie_lo_T28Y84__R2_CONB_0;
  wire tie_lo_T28Y85__R2_CONB_0;
  wire tie_lo_T28Y86__R2_CONB_0;
  wire tie_lo_T28Y87__R2_CONB_0;
  wire tie_lo_T28Y88__R2_CONB_0;
  wire tie_lo_T28Y89__R2_CONB_0;
  wire tie_lo_T28Y8__R2_CONB_0;
  wire tie_lo_T28Y9__R2_CONB_0;
  wire tie_lo_T29Y0__R2_CONB_0;
  wire tie_lo_T29Y10__R2_CONB_0;
  wire tie_lo_T29Y11__R2_CONB_0;
  wire tie_lo_T29Y12__R2_CONB_0;
  wire tie_lo_T29Y13__R2_CONB_0;
  wire tie_lo_T29Y14__R2_CONB_0;
  wire tie_lo_T29Y15__R2_CONB_0;
  wire tie_lo_T29Y16__R2_CONB_0;
  wire tie_lo_T29Y17__R2_CONB_0;
  wire tie_lo_T29Y18__R2_CONB_0;
  wire tie_lo_T29Y19__R2_CONB_0;
  wire tie_lo_T29Y1__R2_CONB_0;
  wire tie_lo_T29Y20__R2_CONB_0;
  wire tie_lo_T29Y21__R2_CONB_0;
  wire tie_lo_T29Y22__R2_CONB_0;
  wire tie_lo_T29Y23__R2_CONB_0;
  wire tie_lo_T29Y24__R2_CONB_0;
  wire tie_lo_T29Y25__R2_CONB_0;
  wire tie_lo_T29Y26__R2_CONB_0;
  wire tie_lo_T29Y27__R2_CONB_0;
  wire tie_lo_T29Y28__R2_CONB_0;
  wire tie_lo_T29Y29__R2_CONB_0;
  wire tie_lo_T29Y2__R2_CONB_0;
  wire tie_lo_T29Y30__R2_CONB_0;
  wire tie_lo_T29Y31__R2_CONB_0;
  wire tie_lo_T29Y32__R2_CONB_0;
  wire tie_lo_T29Y33__R2_CONB_0;
  wire tie_lo_T29Y34__R2_CONB_0;
  wire tie_lo_T29Y35__R2_CONB_0;
  wire tie_lo_T29Y36__R2_CONB_0;
  wire tie_lo_T29Y37__R2_CONB_0;
  wire tie_lo_T29Y38__R2_CONB_0;
  wire tie_lo_T29Y39__R2_CONB_0;
  wire tie_lo_T29Y3__R2_CONB_0;
  wire tie_lo_T29Y40__R2_CONB_0;
  wire tie_lo_T29Y41__R2_CONB_0;
  wire tie_lo_T29Y42__R2_CONB_0;
  wire tie_lo_T29Y43__R2_CONB_0;
  wire tie_lo_T29Y44__R2_CONB_0;
  wire tie_lo_T29Y45__R2_CONB_0;
  wire tie_lo_T29Y46__R2_CONB_0;
  wire tie_lo_T29Y47__R2_CONB_0;
  wire tie_lo_T29Y48__R2_CONB_0;
  wire tie_lo_T29Y49__R2_CONB_0;
  wire tie_lo_T29Y4__R2_CONB_0;
  wire tie_lo_T29Y50__R2_CONB_0;
  wire tie_lo_T29Y51__R2_CONB_0;
  wire tie_lo_T29Y52__R2_CONB_0;
  wire tie_lo_T29Y53__R2_CONB_0;
  wire tie_lo_T29Y54__R2_CONB_0;
  wire tie_lo_T29Y55__R2_CONB_0;
  wire tie_lo_T29Y56__R2_CONB_0;
  wire tie_lo_T29Y57__R2_CONB_0;
  wire tie_lo_T29Y58__R2_CONB_0;
  wire tie_lo_T29Y59__R2_CONB_0;
  wire tie_lo_T29Y5__R2_CONB_0;
  wire tie_lo_T29Y60__R2_CONB_0;
  wire tie_lo_T29Y61__R2_CONB_0;
  wire tie_lo_T29Y62__R2_CONB_0;
  wire tie_lo_T29Y63__R2_CONB_0;
  wire tie_lo_T29Y64__R2_CONB_0;
  wire tie_lo_T29Y65__R2_CONB_0;
  wire tie_lo_T29Y66__R2_CONB_0;
  wire tie_lo_T29Y67__R2_CONB_0;
  wire tie_lo_T29Y68__R2_CONB_0;
  wire tie_lo_T29Y69__R2_CONB_0;
  wire tie_lo_T29Y6__R2_CONB_0;
  wire tie_lo_T29Y70__R2_CONB_0;
  wire tie_lo_T29Y71__R2_CONB_0;
  wire tie_lo_T29Y72__R2_CONB_0;
  wire tie_lo_T29Y73__R2_CONB_0;
  wire tie_lo_T29Y74__R2_CONB_0;
  wire tie_lo_T29Y75__R2_CONB_0;
  wire tie_lo_T29Y76__R2_CONB_0;
  wire tie_lo_T29Y77__R2_CONB_0;
  wire tie_lo_T29Y78__R2_CONB_0;
  wire tie_lo_T29Y79__R2_CONB_0;
  wire tie_lo_T29Y7__R2_CONB_0;
  wire tie_lo_T29Y80__R2_CONB_0;
  wire tie_lo_T29Y81__R2_CONB_0;
  wire tie_lo_T29Y82__R2_CONB_0;
  wire tie_lo_T29Y83__R2_CONB_0;
  wire tie_lo_T29Y84__R2_CONB_0;
  wire tie_lo_T29Y85__R2_CONB_0;
  wire tie_lo_T29Y86__R2_CONB_0;
  wire tie_lo_T29Y87__R2_CONB_0;
  wire tie_lo_T29Y88__R2_CONB_0;
  wire tie_lo_T29Y89__R2_CONB_0;
  wire tie_lo_T29Y8__R2_CONB_0;
  wire tie_lo_T29Y9__R2_CONB_0;
  wire tie_lo_T2Y0__R2_CONB_0;
  wire tie_lo_T2Y10__R2_CONB_0;
  wire tie_lo_T2Y11__R2_CONB_0;
  wire tie_lo_T2Y12__R2_CONB_0;
  wire tie_lo_T2Y13__R2_CONB_0;
  wire tie_lo_T2Y14__R2_CONB_0;
  wire tie_lo_T2Y15__R2_CONB_0;
  wire tie_lo_T2Y16__R2_CONB_0;
  wire tie_lo_T2Y17__R2_CONB_0;
  wire tie_lo_T2Y18__R2_CONB_0;
  wire tie_lo_T2Y19__R2_CONB_0;
  wire tie_lo_T2Y1__R2_CONB_0;
  wire tie_lo_T2Y20__R2_CONB_0;
  wire tie_lo_T2Y21__R2_CONB_0;
  wire tie_lo_T2Y22__R2_CONB_0;
  wire tie_lo_T2Y23__R2_CONB_0;
  wire tie_lo_T2Y24__R2_CONB_0;
  wire tie_lo_T2Y25__R2_CONB_0;
  wire tie_lo_T2Y26__R2_CONB_0;
  wire tie_lo_T2Y27__R2_CONB_0;
  wire tie_lo_T2Y28__R2_CONB_0;
  wire tie_lo_T2Y29__R2_CONB_0;
  wire tie_lo_T2Y2__R2_CONB_0;
  wire tie_lo_T2Y30__R2_CONB_0;
  wire tie_lo_T2Y31__R2_CONB_0;
  wire tie_lo_T2Y32__R2_CONB_0;
  wire tie_lo_T2Y33__R2_CONB_0;
  wire tie_lo_T2Y34__R2_CONB_0;
  wire tie_lo_T2Y35__R2_CONB_0;
  wire tie_lo_T2Y36__R2_CONB_0;
  wire tie_lo_T2Y37__R2_CONB_0;
  wire tie_lo_T2Y38__R2_CONB_0;
  wire tie_lo_T2Y39__R2_CONB_0;
  wire tie_lo_T2Y3__R2_CONB_0;
  wire tie_lo_T2Y40__R2_CONB_0;
  wire tie_lo_T2Y41__R2_CONB_0;
  wire tie_lo_T2Y42__R2_CONB_0;
  wire tie_lo_T2Y43__R2_CONB_0;
  wire tie_lo_T2Y44__R2_CONB_0;
  wire tie_lo_T2Y45__R2_CONB_0;
  wire tie_lo_T2Y46__R2_CONB_0;
  wire tie_lo_T2Y47__R2_CONB_0;
  wire tie_lo_T2Y48__R2_CONB_0;
  wire tie_lo_T2Y49__R2_CONB_0;
  wire tie_lo_T2Y4__R2_CONB_0;
  wire tie_lo_T2Y50__R2_CONB_0;
  wire tie_lo_T2Y51__R2_CONB_0;
  wire tie_lo_T2Y52__R2_CONB_0;
  wire tie_lo_T2Y53__R2_CONB_0;
  wire tie_lo_T2Y54__R2_CONB_0;
  wire tie_lo_T2Y55__R2_CONB_0;
  wire tie_lo_T2Y56__R2_CONB_0;
  wire tie_lo_T2Y57__R2_CONB_0;
  wire tie_lo_T2Y58__R2_CONB_0;
  wire tie_lo_T2Y59__R2_CONB_0;
  wire tie_lo_T2Y5__R2_CONB_0;
  wire tie_lo_T2Y60__R2_CONB_0;
  wire tie_lo_T2Y61__R2_CONB_0;
  wire tie_lo_T2Y62__R2_CONB_0;
  wire tie_lo_T2Y63__R2_CONB_0;
  wire tie_lo_T2Y64__R2_CONB_0;
  wire tie_lo_T2Y65__R2_CONB_0;
  wire tie_lo_T2Y66__R2_CONB_0;
  wire tie_lo_T2Y67__R2_CONB_0;
  wire tie_lo_T2Y68__R2_CONB_0;
  wire tie_lo_T2Y69__R2_CONB_0;
  wire tie_lo_T2Y6__R2_CONB_0;
  wire tie_lo_T2Y70__R2_CONB_0;
  wire tie_lo_T2Y71__R2_CONB_0;
  wire tie_lo_T2Y72__R2_CONB_0;
  wire tie_lo_T2Y73__R2_CONB_0;
  wire tie_lo_T2Y74__R2_CONB_0;
  wire tie_lo_T2Y75__R2_CONB_0;
  wire tie_lo_T2Y76__R2_CONB_0;
  wire tie_lo_T2Y77__R2_CONB_0;
  wire tie_lo_T2Y78__R2_CONB_0;
  wire tie_lo_T2Y79__R2_CONB_0;
  wire tie_lo_T2Y7__R2_CONB_0;
  wire tie_lo_T2Y80__R2_CONB_0;
  wire tie_lo_T2Y81__R2_CONB_0;
  wire tie_lo_T2Y82__R2_CONB_0;
  wire tie_lo_T2Y83__R2_CONB_0;
  wire tie_lo_T2Y84__R2_CONB_0;
  wire tie_lo_T2Y85__R2_CONB_0;
  wire tie_lo_T2Y86__R2_CONB_0;
  wire tie_lo_T2Y87__R2_CONB_0;
  wire tie_lo_T2Y88__R2_CONB_0;
  wire tie_lo_T2Y89__R2_CONB_0;
  wire tie_lo_T2Y8__R2_CONB_0;
  wire tie_lo_T2Y9__R2_CONB_0;
  wire tie_lo_T30Y0__R2_CONB_0;
  wire tie_lo_T30Y10__R2_CONB_0;
  wire tie_lo_T30Y11__R2_CONB_0;
  wire tie_lo_T30Y12__R2_CONB_0;
  wire tie_lo_T30Y13__R2_CONB_0;
  wire tie_lo_T30Y14__R2_CONB_0;
  wire tie_lo_T30Y15__R2_CONB_0;
  wire tie_lo_T30Y16__R2_CONB_0;
  wire tie_lo_T30Y17__R2_CONB_0;
  wire tie_lo_T30Y18__R2_CONB_0;
  wire tie_lo_T30Y19__R2_CONB_0;
  wire tie_lo_T30Y1__R2_CONB_0;
  wire tie_lo_T30Y20__R2_CONB_0;
  wire tie_lo_T30Y21__R2_CONB_0;
  wire tie_lo_T30Y22__R2_CONB_0;
  wire tie_lo_T30Y23__R2_CONB_0;
  wire tie_lo_T30Y24__R2_CONB_0;
  wire tie_lo_T30Y25__R2_CONB_0;
  wire tie_lo_T30Y26__R2_CONB_0;
  wire tie_lo_T30Y27__R2_CONB_0;
  wire tie_lo_T30Y28__R2_CONB_0;
  wire tie_lo_T30Y29__R2_CONB_0;
  wire tie_lo_T30Y2__R2_CONB_0;
  wire tie_lo_T30Y30__R2_CONB_0;
  wire tie_lo_T30Y31__R2_CONB_0;
  wire tie_lo_T30Y32__R2_CONB_0;
  wire tie_lo_T30Y33__R2_CONB_0;
  wire tie_lo_T30Y34__R2_CONB_0;
  wire tie_lo_T30Y35__R2_CONB_0;
  wire tie_lo_T30Y36__R2_CONB_0;
  wire tie_lo_T30Y37__R2_CONB_0;
  wire tie_lo_T30Y38__R2_CONB_0;
  wire tie_lo_T30Y39__R2_CONB_0;
  wire tie_lo_T30Y3__R2_CONB_0;
  wire tie_lo_T30Y40__R2_CONB_0;
  wire tie_lo_T30Y41__R2_CONB_0;
  wire tie_lo_T30Y42__R2_CONB_0;
  wire tie_lo_T30Y43__R2_CONB_0;
  wire tie_lo_T30Y44__R2_CONB_0;
  wire tie_lo_T30Y45__R2_CONB_0;
  wire tie_lo_T30Y46__R2_CONB_0;
  wire tie_lo_T30Y47__R2_CONB_0;
  wire tie_lo_T30Y48__R2_CONB_0;
  wire tie_lo_T30Y49__R2_CONB_0;
  wire tie_lo_T30Y4__R2_CONB_0;
  wire tie_lo_T30Y50__R2_CONB_0;
  wire tie_lo_T30Y51__R2_CONB_0;
  wire tie_lo_T30Y52__R2_CONB_0;
  wire tie_lo_T30Y53__R2_CONB_0;
  wire tie_lo_T30Y54__R2_CONB_0;
  wire tie_lo_T30Y55__R2_CONB_0;
  wire tie_lo_T30Y56__R2_CONB_0;
  wire tie_lo_T30Y57__R2_CONB_0;
  wire tie_lo_T30Y58__R2_CONB_0;
  wire tie_lo_T30Y59__R2_CONB_0;
  wire tie_lo_T30Y5__R2_CONB_0;
  wire tie_lo_T30Y60__R2_CONB_0;
  wire tie_lo_T30Y61__R2_CONB_0;
  wire tie_lo_T30Y62__R2_CONB_0;
  wire tie_lo_T30Y63__R2_CONB_0;
  wire tie_lo_T30Y64__R2_CONB_0;
  wire tie_lo_T30Y65__R2_CONB_0;
  wire tie_lo_T30Y66__R2_CONB_0;
  wire tie_lo_T30Y67__R2_CONB_0;
  wire tie_lo_T30Y68__R2_CONB_0;
  wire tie_lo_T30Y69__R2_CONB_0;
  wire tie_lo_T30Y6__R2_CONB_0;
  wire tie_lo_T30Y70__R2_CONB_0;
  wire tie_lo_T30Y71__R2_CONB_0;
  wire tie_lo_T30Y72__R2_CONB_0;
  wire tie_lo_T30Y73__R2_CONB_0;
  wire tie_lo_T30Y74__R2_CONB_0;
  wire tie_lo_T30Y75__R2_CONB_0;
  wire tie_lo_T30Y76__R2_CONB_0;
  wire tie_lo_T30Y77__R2_CONB_0;
  wire tie_lo_T30Y78__R2_CONB_0;
  wire tie_lo_T30Y79__R2_CONB_0;
  wire tie_lo_T30Y7__R2_CONB_0;
  wire tie_lo_T30Y80__R2_CONB_0;
  wire tie_lo_T30Y81__R2_CONB_0;
  wire tie_lo_T30Y82__R2_CONB_0;
  wire tie_lo_T30Y83__R2_CONB_0;
  wire tie_lo_T30Y84__R2_CONB_0;
  wire tie_lo_T30Y85__R2_CONB_0;
  wire tie_lo_T30Y86__R2_CONB_0;
  wire tie_lo_T30Y87__R2_CONB_0;
  wire tie_lo_T30Y88__R2_CONB_0;
  wire tie_lo_T30Y89__R2_CONB_0;
  wire tie_lo_T30Y8__R2_CONB_0;
  wire tie_lo_T30Y9__R2_CONB_0;
  wire tie_lo_T31Y0__R2_CONB_0;
  wire tie_lo_T31Y10__R2_CONB_0;
  wire tie_lo_T31Y11__R2_CONB_0;
  wire tie_lo_T31Y12__R2_CONB_0;
  wire tie_lo_T31Y13__R2_CONB_0;
  wire tie_lo_T31Y14__R2_CONB_0;
  wire tie_lo_T31Y15__R2_CONB_0;
  wire tie_lo_T31Y16__R2_CONB_0;
  wire tie_lo_T31Y17__R2_CONB_0;
  wire tie_lo_T31Y18__R2_CONB_0;
  wire tie_lo_T31Y19__R2_CONB_0;
  wire tie_lo_T31Y1__R2_CONB_0;
  wire tie_lo_T31Y20__R2_CONB_0;
  wire tie_lo_T31Y21__R2_CONB_0;
  wire tie_lo_T31Y22__R2_CONB_0;
  wire tie_lo_T31Y23__R2_CONB_0;
  wire tie_lo_T31Y24__R2_CONB_0;
  wire tie_lo_T31Y25__R2_CONB_0;
  wire tie_lo_T31Y26__R2_CONB_0;
  wire tie_lo_T31Y27__R2_CONB_0;
  wire tie_lo_T31Y28__R2_CONB_0;
  wire tie_lo_T31Y29__R2_CONB_0;
  wire tie_lo_T31Y2__R2_CONB_0;
  wire tie_lo_T31Y30__R2_CONB_0;
  wire tie_lo_T31Y31__R2_CONB_0;
  wire tie_lo_T31Y32__R2_CONB_0;
  wire tie_lo_T31Y33__R2_CONB_0;
  wire tie_lo_T31Y34__R2_CONB_0;
  wire tie_lo_T31Y35__R2_CONB_0;
  wire tie_lo_T31Y36__R2_CONB_0;
  wire tie_lo_T31Y37__R2_CONB_0;
  wire tie_lo_T31Y38__R2_CONB_0;
  wire tie_lo_T31Y39__R2_CONB_0;
  wire tie_lo_T31Y3__R2_CONB_0;
  wire tie_lo_T31Y40__R2_CONB_0;
  wire tie_lo_T31Y41__R2_CONB_0;
  wire tie_lo_T31Y42__R2_CONB_0;
  wire tie_lo_T31Y43__R2_CONB_0;
  wire tie_lo_T31Y44__R2_CONB_0;
  wire tie_lo_T31Y45__R2_CONB_0;
  wire tie_lo_T31Y46__R2_CONB_0;
  wire tie_lo_T31Y47__R2_CONB_0;
  wire tie_lo_T31Y48__R2_CONB_0;
  wire tie_lo_T31Y49__R2_CONB_0;
  wire tie_lo_T31Y4__R2_CONB_0;
  wire tie_lo_T31Y50__R2_CONB_0;
  wire tie_lo_T31Y51__R2_CONB_0;
  wire tie_lo_T31Y52__R2_CONB_0;
  wire tie_lo_T31Y53__R2_CONB_0;
  wire tie_lo_T31Y54__R2_CONB_0;
  wire tie_lo_T31Y55__R2_CONB_0;
  wire tie_lo_T31Y56__R2_CONB_0;
  wire tie_lo_T31Y57__R2_CONB_0;
  wire tie_lo_T31Y58__R2_CONB_0;
  wire tie_lo_T31Y59__R2_CONB_0;
  wire tie_lo_T31Y5__R2_CONB_0;
  wire tie_lo_T31Y60__R2_CONB_0;
  wire tie_lo_T31Y61__R2_CONB_0;
  wire tie_lo_T31Y62__R2_CONB_0;
  wire tie_lo_T31Y63__R2_CONB_0;
  wire tie_lo_T31Y64__R2_CONB_0;
  wire tie_lo_T31Y65__R2_CONB_0;
  wire tie_lo_T31Y66__R2_CONB_0;
  wire tie_lo_T31Y67__R2_CONB_0;
  wire tie_lo_T31Y68__R2_CONB_0;
  wire tie_lo_T31Y69__R2_CONB_0;
  wire tie_lo_T31Y6__R2_CONB_0;
  wire tie_lo_T31Y70__R2_CONB_0;
  wire tie_lo_T31Y71__R2_CONB_0;
  wire tie_lo_T31Y72__R2_CONB_0;
  wire tie_lo_T31Y73__R2_CONB_0;
  wire tie_lo_T31Y74__R2_CONB_0;
  wire tie_lo_T31Y75__R2_CONB_0;
  wire tie_lo_T31Y76__R2_CONB_0;
  wire tie_lo_T31Y77__R2_CONB_0;
  wire tie_lo_T31Y78__R2_CONB_0;
  wire tie_lo_T31Y79__R2_CONB_0;
  wire tie_lo_T31Y7__R2_CONB_0;
  wire tie_lo_T31Y80__R2_CONB_0;
  wire tie_lo_T31Y81__R2_CONB_0;
  wire tie_lo_T31Y82__R2_CONB_0;
  wire tie_lo_T31Y83__R2_CONB_0;
  wire tie_lo_T31Y84__R2_CONB_0;
  wire tie_lo_T31Y85__R2_CONB_0;
  wire tie_lo_T31Y86__R2_CONB_0;
  wire tie_lo_T31Y87__R2_CONB_0;
  wire tie_lo_T31Y88__R2_CONB_0;
  wire tie_lo_T31Y89__R2_CONB_0;
  wire tie_lo_T31Y8__R2_CONB_0;
  wire tie_lo_T31Y9__R2_CONB_0;
  wire tie_lo_T32Y0__R2_CONB_0;
  wire tie_lo_T32Y10__R2_CONB_0;
  wire tie_lo_T32Y11__R2_CONB_0;
  wire tie_lo_T32Y12__R2_CONB_0;
  wire tie_lo_T32Y13__R2_CONB_0;
  wire tie_lo_T32Y14__R2_CONB_0;
  wire tie_lo_T32Y15__R2_CONB_0;
  wire tie_lo_T32Y16__R2_CONB_0;
  wire tie_lo_T32Y17__R2_CONB_0;
  wire tie_lo_T32Y18__R2_CONB_0;
  wire tie_lo_T32Y19__R2_CONB_0;
  wire tie_lo_T32Y1__R2_CONB_0;
  wire tie_lo_T32Y20__R2_CONB_0;
  wire tie_lo_T32Y21__R2_CONB_0;
  wire tie_lo_T32Y22__R2_CONB_0;
  wire tie_lo_T32Y23__R2_CONB_0;
  wire tie_lo_T32Y24__R2_CONB_0;
  wire tie_lo_T32Y25__R2_CONB_0;
  wire tie_lo_T32Y26__R2_CONB_0;
  wire tie_lo_T32Y27__R2_CONB_0;
  wire tie_lo_T32Y28__R2_CONB_0;
  wire tie_lo_T32Y29__R2_CONB_0;
  wire tie_lo_T32Y2__R2_CONB_0;
  wire tie_lo_T32Y30__R2_CONB_0;
  wire tie_lo_T32Y31__R2_CONB_0;
  wire tie_lo_T32Y32__R2_CONB_0;
  wire tie_lo_T32Y33__R2_CONB_0;
  wire tie_lo_T32Y34__R2_CONB_0;
  wire tie_lo_T32Y35__R2_CONB_0;
  wire tie_lo_T32Y36__R2_CONB_0;
  wire tie_lo_T32Y37__R2_CONB_0;
  wire tie_lo_T32Y38__R2_CONB_0;
  wire tie_lo_T32Y39__R2_CONB_0;
  wire tie_lo_T32Y3__R2_CONB_0;
  wire tie_lo_T32Y40__R2_CONB_0;
  wire tie_lo_T32Y41__R2_CONB_0;
  wire tie_lo_T32Y42__R2_CONB_0;
  wire tie_lo_T32Y43__R2_CONB_0;
  wire tie_lo_T32Y44__R2_CONB_0;
  wire tie_lo_T32Y45__R2_CONB_0;
  wire tie_lo_T32Y46__R2_CONB_0;
  wire tie_lo_T32Y47__R2_CONB_0;
  wire tie_lo_T32Y48__R2_CONB_0;
  wire tie_lo_T32Y49__R2_CONB_0;
  wire tie_lo_T32Y4__R2_CONB_0;
  wire tie_lo_T32Y50__R2_CONB_0;
  wire tie_lo_T32Y51__R2_CONB_0;
  wire tie_lo_T32Y52__R2_CONB_0;
  wire tie_lo_T32Y53__R2_CONB_0;
  wire tie_lo_T32Y54__R2_CONB_0;
  wire tie_lo_T32Y55__R2_CONB_0;
  wire tie_lo_T32Y56__R2_CONB_0;
  wire tie_lo_T32Y57__R2_CONB_0;
  wire tie_lo_T32Y58__R2_CONB_0;
  wire tie_lo_T32Y59__R2_CONB_0;
  wire tie_lo_T32Y5__R2_CONB_0;
  wire tie_lo_T32Y60__R2_CONB_0;
  wire tie_lo_T32Y61__R2_CONB_0;
  wire tie_lo_T32Y62__R2_CONB_0;
  wire tie_lo_T32Y63__R2_CONB_0;
  wire tie_lo_T32Y64__R2_CONB_0;
  wire tie_lo_T32Y65__R2_CONB_0;
  wire tie_lo_T32Y66__R2_CONB_0;
  wire tie_lo_T32Y67__R2_CONB_0;
  wire tie_lo_T32Y68__R2_CONB_0;
  wire tie_lo_T32Y69__R2_CONB_0;
  wire tie_lo_T32Y6__R2_CONB_0;
  wire tie_lo_T32Y70__R2_CONB_0;
  wire tie_lo_T32Y71__R2_CONB_0;
  wire tie_lo_T32Y72__R2_CONB_0;
  wire tie_lo_T32Y73__R2_CONB_0;
  wire tie_lo_T32Y74__R2_CONB_0;
  wire tie_lo_T32Y75__R2_CONB_0;
  wire tie_lo_T32Y76__R2_CONB_0;
  wire tie_lo_T32Y77__R2_CONB_0;
  wire tie_lo_T32Y78__R2_CONB_0;
  wire tie_lo_T32Y79__R2_CONB_0;
  wire tie_lo_T32Y7__R2_CONB_0;
  wire tie_lo_T32Y80__R2_CONB_0;
  wire tie_lo_T32Y81__R2_CONB_0;
  wire tie_lo_T32Y82__R2_CONB_0;
  wire tie_lo_T32Y83__R2_CONB_0;
  wire tie_lo_T32Y84__R2_CONB_0;
  wire tie_lo_T32Y85__R2_CONB_0;
  wire tie_lo_T32Y86__R2_CONB_0;
  wire tie_lo_T32Y87__R2_CONB_0;
  wire tie_lo_T32Y88__R2_CONB_0;
  wire tie_lo_T32Y89__R2_CONB_0;
  wire tie_lo_T32Y8__R2_CONB_0;
  wire tie_lo_T32Y9__R2_CONB_0;
  wire tie_lo_T33Y0__R2_CONB_0;
  wire tie_lo_T33Y10__R2_CONB_0;
  wire tie_lo_T33Y11__R2_CONB_0;
  wire tie_lo_T33Y12__R2_CONB_0;
  wire tie_lo_T33Y13__R2_CONB_0;
  wire tie_lo_T33Y14__R2_CONB_0;
  wire tie_lo_T33Y15__R2_CONB_0;
  wire tie_lo_T33Y16__R2_CONB_0;
  wire tie_lo_T33Y17__R2_CONB_0;
  wire tie_lo_T33Y18__R2_CONB_0;
  wire tie_lo_T33Y19__R2_CONB_0;
  wire tie_lo_T33Y1__R2_CONB_0;
  wire tie_lo_T33Y20__R2_CONB_0;
  wire tie_lo_T33Y21__R2_CONB_0;
  wire tie_lo_T33Y22__R2_CONB_0;
  wire tie_lo_T33Y23__R2_CONB_0;
  wire tie_lo_T33Y24__R2_CONB_0;
  wire tie_lo_T33Y25__R2_CONB_0;
  wire tie_lo_T33Y26__R2_CONB_0;
  wire tie_lo_T33Y27__R2_CONB_0;
  wire tie_lo_T33Y28__R2_CONB_0;
  wire tie_lo_T33Y29__R2_CONB_0;
  wire tie_lo_T33Y2__R2_CONB_0;
  wire tie_lo_T33Y30__R2_CONB_0;
  wire tie_lo_T33Y31__R2_CONB_0;
  wire tie_lo_T33Y32__R2_CONB_0;
  wire tie_lo_T33Y33__R2_CONB_0;
  wire tie_lo_T33Y34__R2_CONB_0;
  wire tie_lo_T33Y35__R2_CONB_0;
  wire tie_lo_T33Y36__R2_CONB_0;
  wire tie_lo_T33Y37__R2_CONB_0;
  wire tie_lo_T33Y38__R2_CONB_0;
  wire tie_lo_T33Y39__R2_CONB_0;
  wire tie_lo_T33Y3__R2_CONB_0;
  wire tie_lo_T33Y40__R2_CONB_0;
  wire tie_lo_T33Y41__R2_CONB_0;
  wire tie_lo_T33Y42__R2_CONB_0;
  wire tie_lo_T33Y43__R2_CONB_0;
  wire tie_lo_T33Y44__R2_CONB_0;
  wire tie_lo_T33Y45__R2_CONB_0;
  wire tie_lo_T33Y46__R2_CONB_0;
  wire tie_lo_T33Y47__R2_CONB_0;
  wire tie_lo_T33Y48__R2_CONB_0;
  wire tie_lo_T33Y49__R2_CONB_0;
  wire tie_lo_T33Y4__R2_CONB_0;
  wire tie_lo_T33Y50__R2_CONB_0;
  wire tie_lo_T33Y51__R2_CONB_0;
  wire tie_lo_T33Y52__R2_CONB_0;
  wire tie_lo_T33Y53__R2_CONB_0;
  wire tie_lo_T33Y54__R2_CONB_0;
  wire tie_lo_T33Y55__R2_CONB_0;
  wire tie_lo_T33Y56__R2_CONB_0;
  wire tie_lo_T33Y57__R2_CONB_0;
  wire tie_lo_T33Y58__R2_CONB_0;
  wire tie_lo_T33Y59__R2_CONB_0;
  wire tie_lo_T33Y5__R2_CONB_0;
  wire tie_lo_T33Y60__R2_CONB_0;
  wire tie_lo_T33Y61__R2_CONB_0;
  wire tie_lo_T33Y62__R2_CONB_0;
  wire tie_lo_T33Y63__R2_CONB_0;
  wire tie_lo_T33Y64__R2_CONB_0;
  wire tie_lo_T33Y65__R2_CONB_0;
  wire tie_lo_T33Y66__R2_CONB_0;
  wire tie_lo_T33Y67__R2_CONB_0;
  wire tie_lo_T33Y68__R2_CONB_0;
  wire tie_lo_T33Y69__R2_CONB_0;
  wire tie_lo_T33Y6__R2_CONB_0;
  wire tie_lo_T33Y70__R2_CONB_0;
  wire tie_lo_T33Y71__R2_CONB_0;
  wire tie_lo_T33Y72__R2_CONB_0;
  wire tie_lo_T33Y73__R2_CONB_0;
  wire tie_lo_T33Y74__R2_CONB_0;
  wire tie_lo_T33Y75__R2_CONB_0;
  wire tie_lo_T33Y76__R2_CONB_0;
  wire tie_lo_T33Y77__R2_CONB_0;
  wire tie_lo_T33Y78__R2_CONB_0;
  wire tie_lo_T33Y79__R2_CONB_0;
  wire tie_lo_T33Y7__R2_CONB_0;
  wire tie_lo_T33Y80__R2_CONB_0;
  wire tie_lo_T33Y81__R2_CONB_0;
  wire tie_lo_T33Y82__R2_CONB_0;
  wire tie_lo_T33Y83__R2_CONB_0;
  wire tie_lo_T33Y84__R2_CONB_0;
  wire tie_lo_T33Y85__R2_CONB_0;
  wire tie_lo_T33Y86__R2_CONB_0;
  wire tie_lo_T33Y87__R2_CONB_0;
  wire tie_lo_T33Y88__R2_CONB_0;
  wire tie_lo_T33Y89__R2_CONB_0;
  wire tie_lo_T33Y8__R2_CONB_0;
  wire tie_lo_T33Y9__R2_CONB_0;
  wire tie_lo_T34Y0__R2_CONB_0;
  wire tie_lo_T34Y10__R2_CONB_0;
  wire tie_lo_T34Y11__R2_CONB_0;
  wire tie_lo_T34Y12__R2_CONB_0;
  wire tie_lo_T34Y13__R2_CONB_0;
  wire tie_lo_T34Y14__R2_CONB_0;
  wire tie_lo_T34Y15__R2_CONB_0;
  wire tie_lo_T34Y16__R2_CONB_0;
  wire tie_lo_T34Y17__R2_CONB_0;
  wire tie_lo_T34Y18__R2_CONB_0;
  wire tie_lo_T34Y19__R2_CONB_0;
  wire tie_lo_T34Y1__R2_CONB_0;
  wire tie_lo_T34Y20__R2_CONB_0;
  wire tie_lo_T34Y21__R2_CONB_0;
  wire tie_lo_T34Y22__R2_CONB_0;
  wire tie_lo_T34Y23__R2_CONB_0;
  wire tie_lo_T34Y24__R2_CONB_0;
  wire tie_lo_T34Y25__R2_CONB_0;
  wire tie_lo_T34Y26__R2_CONB_0;
  wire tie_lo_T34Y27__R2_CONB_0;
  wire tie_lo_T34Y28__R2_CONB_0;
  wire tie_lo_T34Y29__R2_CONB_0;
  wire tie_lo_T34Y2__R2_CONB_0;
  wire tie_lo_T34Y30__R2_CONB_0;
  wire tie_lo_T34Y31__R2_CONB_0;
  wire tie_lo_T34Y32__R2_CONB_0;
  wire tie_lo_T34Y33__R2_CONB_0;
  wire tie_lo_T34Y34__R2_CONB_0;
  wire tie_lo_T34Y35__R2_CONB_0;
  wire tie_lo_T34Y36__R2_CONB_0;
  wire tie_lo_T34Y37__R2_CONB_0;
  wire tie_lo_T34Y38__R2_CONB_0;
  wire tie_lo_T34Y39__R2_CONB_0;
  wire tie_lo_T34Y3__R2_CONB_0;
  wire tie_lo_T34Y40__R2_CONB_0;
  wire tie_lo_T34Y41__R2_CONB_0;
  wire tie_lo_T34Y42__R2_CONB_0;
  wire tie_lo_T34Y43__R2_CONB_0;
  wire tie_lo_T34Y44__R2_CONB_0;
  wire tie_lo_T34Y45__R2_CONB_0;
  wire tie_lo_T34Y46__R2_CONB_0;
  wire tie_lo_T34Y47__R2_CONB_0;
  wire tie_lo_T34Y48__R2_CONB_0;
  wire tie_lo_T34Y49__R2_CONB_0;
  wire tie_lo_T34Y4__R2_CONB_0;
  wire tie_lo_T34Y50__R2_CONB_0;
  wire tie_lo_T34Y51__R2_CONB_0;
  wire tie_lo_T34Y52__R2_CONB_0;
  wire tie_lo_T34Y53__R2_CONB_0;
  wire tie_lo_T34Y54__R2_CONB_0;
  wire tie_lo_T34Y55__R2_CONB_0;
  wire tie_lo_T34Y56__R2_CONB_0;
  wire tie_lo_T34Y57__R2_CONB_0;
  wire tie_lo_T34Y58__R2_CONB_0;
  wire tie_lo_T34Y59__R2_CONB_0;
  wire tie_lo_T34Y5__R2_CONB_0;
  wire tie_lo_T34Y60__R2_CONB_0;
  wire tie_lo_T34Y61__R2_CONB_0;
  wire tie_lo_T34Y62__R2_CONB_0;
  wire tie_lo_T34Y63__R2_CONB_0;
  wire tie_lo_T34Y64__R2_CONB_0;
  wire tie_lo_T34Y65__R2_CONB_0;
  wire tie_lo_T34Y66__R2_CONB_0;
  wire tie_lo_T34Y67__R2_CONB_0;
  wire tie_lo_T34Y68__R2_CONB_0;
  wire tie_lo_T34Y69__R2_CONB_0;
  wire tie_lo_T34Y6__R2_CONB_0;
  wire tie_lo_T34Y70__R2_CONB_0;
  wire tie_lo_T34Y71__R2_CONB_0;
  wire tie_lo_T34Y72__R2_CONB_0;
  wire tie_lo_T34Y73__R2_CONB_0;
  wire tie_lo_T34Y74__R2_CONB_0;
  wire tie_lo_T34Y75__R2_CONB_0;
  wire tie_lo_T34Y76__R2_CONB_0;
  wire tie_lo_T34Y77__R2_CONB_0;
  wire tie_lo_T34Y78__R2_CONB_0;
  wire tie_lo_T34Y79__R2_CONB_0;
  wire tie_lo_T34Y7__R2_CONB_0;
  wire tie_lo_T34Y80__R2_CONB_0;
  wire tie_lo_T34Y81__R2_CONB_0;
  wire tie_lo_T34Y82__R2_CONB_0;
  wire tie_lo_T34Y83__R2_CONB_0;
  wire tie_lo_T34Y84__R2_CONB_0;
  wire tie_lo_T34Y85__R2_CONB_0;
  wire tie_lo_T34Y86__R2_CONB_0;
  wire tie_lo_T34Y87__R2_CONB_0;
  wire tie_lo_T34Y88__R2_CONB_0;
  wire tie_lo_T34Y89__R2_CONB_0;
  wire tie_lo_T34Y8__R2_CONB_0;
  wire tie_lo_T34Y9__R2_CONB_0;
  wire tie_lo_T35Y0__R2_CONB_0;
  wire tie_lo_T35Y10__R2_CONB_0;
  wire tie_lo_T35Y11__R2_CONB_0;
  wire tie_lo_T35Y12__R2_CONB_0;
  wire tie_lo_T35Y13__R2_CONB_0;
  wire tie_lo_T35Y14__R2_CONB_0;
  wire tie_lo_T35Y15__R2_CONB_0;
  wire tie_lo_T35Y16__R2_CONB_0;
  wire tie_lo_T35Y17__R2_CONB_0;
  wire tie_lo_T35Y18__R2_CONB_0;
  wire tie_lo_T35Y19__R2_CONB_0;
  wire tie_lo_T35Y1__R2_CONB_0;
  wire tie_lo_T35Y20__R2_CONB_0;
  wire tie_lo_T35Y21__R2_CONB_0;
  wire tie_lo_T35Y22__R2_CONB_0;
  wire tie_lo_T35Y23__R2_CONB_0;
  wire tie_lo_T35Y24__R2_CONB_0;
  wire tie_lo_T35Y25__R2_CONB_0;
  wire tie_lo_T35Y26__R2_CONB_0;
  wire tie_lo_T35Y27__R2_CONB_0;
  wire tie_lo_T35Y28__R2_CONB_0;
  wire tie_lo_T35Y29__R2_CONB_0;
  wire tie_lo_T35Y2__R2_CONB_0;
  wire tie_lo_T35Y30__R2_CONB_0;
  wire tie_lo_T35Y31__R2_CONB_0;
  wire tie_lo_T35Y32__R2_CONB_0;
  wire tie_lo_T35Y33__R2_CONB_0;
  wire tie_lo_T35Y34__R2_CONB_0;
  wire tie_lo_T35Y35__R2_CONB_0;
  wire tie_lo_T35Y36__R2_CONB_0;
  wire tie_lo_T35Y37__R2_CONB_0;
  wire tie_lo_T35Y38__R2_CONB_0;
  wire tie_lo_T35Y39__R2_CONB_0;
  wire tie_lo_T35Y3__R2_CONB_0;
  wire tie_lo_T35Y40__R2_CONB_0;
  wire tie_lo_T35Y41__R2_CONB_0;
  wire tie_lo_T35Y42__R2_CONB_0;
  wire tie_lo_T35Y43__R2_CONB_0;
  wire tie_lo_T35Y44__R2_CONB_0;
  wire tie_lo_T35Y45__R2_CONB_0;
  wire tie_lo_T35Y46__R2_CONB_0;
  wire tie_lo_T35Y47__R2_CONB_0;
  wire tie_lo_T35Y48__R2_CONB_0;
  wire tie_lo_T35Y49__R2_CONB_0;
  wire tie_lo_T35Y4__R2_CONB_0;
  wire tie_lo_T35Y50__R2_CONB_0;
  wire tie_lo_T35Y51__R2_CONB_0;
  wire tie_lo_T35Y52__R2_CONB_0;
  wire tie_lo_T35Y53__R2_CONB_0;
  wire tie_lo_T35Y54__R2_CONB_0;
  wire tie_lo_T35Y55__R2_CONB_0;
  wire tie_lo_T35Y56__R2_CONB_0;
  wire tie_lo_T35Y57__R2_CONB_0;
  wire tie_lo_T35Y58__R2_CONB_0;
  wire tie_lo_T35Y59__R2_CONB_0;
  wire tie_lo_T35Y5__R2_CONB_0;
  wire tie_lo_T35Y60__R2_CONB_0;
  wire tie_lo_T35Y61__R2_CONB_0;
  wire tie_lo_T35Y62__R2_CONB_0;
  wire tie_lo_T35Y63__R2_CONB_0;
  wire tie_lo_T35Y64__R2_CONB_0;
  wire tie_lo_T35Y65__R2_CONB_0;
  wire tie_lo_T35Y66__R2_CONB_0;
  wire tie_lo_T35Y67__R2_CONB_0;
  wire tie_lo_T35Y68__R2_CONB_0;
  wire tie_lo_T35Y69__R2_CONB_0;
  wire tie_lo_T35Y6__R2_CONB_0;
  wire tie_lo_T35Y70__R2_CONB_0;
  wire tie_lo_T35Y71__R2_CONB_0;
  wire tie_lo_T35Y72__R2_CONB_0;
  wire tie_lo_T35Y73__R2_CONB_0;
  wire tie_lo_T35Y74__R2_CONB_0;
  wire tie_lo_T35Y75__R2_CONB_0;
  wire tie_lo_T35Y76__R2_CONB_0;
  wire tie_lo_T35Y77__R2_CONB_0;
  wire tie_lo_T35Y78__R2_CONB_0;
  wire tie_lo_T35Y79__R2_CONB_0;
  wire tie_lo_T35Y7__R2_CONB_0;
  wire tie_lo_T35Y80__R2_CONB_0;
  wire tie_lo_T35Y81__R2_CONB_0;
  wire tie_lo_T35Y82__R2_CONB_0;
  wire tie_lo_T35Y83__R2_CONB_0;
  wire tie_lo_T35Y84__R2_CONB_0;
  wire tie_lo_T35Y85__R2_CONB_0;
  wire tie_lo_T35Y86__R2_CONB_0;
  wire tie_lo_T35Y87__R2_CONB_0;
  wire tie_lo_T35Y88__R2_CONB_0;
  wire tie_lo_T35Y89__R2_CONB_0;
  wire tie_lo_T35Y8__R2_CONB_0;
  wire tie_lo_T35Y9__R2_CONB_0;
  wire tie_lo_T3Y0__R2_CONB_0;
  wire tie_lo_T3Y10__R2_CONB_0;
  wire tie_lo_T3Y11__R2_CONB_0;
  wire tie_lo_T3Y12__R2_CONB_0;
  wire tie_lo_T3Y13__R2_CONB_0;
  wire tie_lo_T3Y14__R2_CONB_0;
  wire tie_lo_T3Y15__R2_CONB_0;
  wire tie_lo_T3Y16__R2_CONB_0;
  wire tie_lo_T3Y17__R2_CONB_0;
  wire tie_lo_T3Y18__R2_CONB_0;
  wire tie_lo_T3Y19__R2_CONB_0;
  wire tie_lo_T3Y1__R2_CONB_0;
  wire tie_lo_T3Y20__R2_CONB_0;
  wire tie_lo_T3Y21__R2_CONB_0;
  wire tie_lo_T3Y22__R2_CONB_0;
  wire tie_lo_T3Y23__R2_CONB_0;
  wire tie_lo_T3Y24__R2_CONB_0;
  wire tie_lo_T3Y25__R2_CONB_0;
  wire tie_lo_T3Y26__R2_CONB_0;
  wire tie_lo_T3Y27__R2_CONB_0;
  wire tie_lo_T3Y28__R2_CONB_0;
  wire tie_lo_T3Y29__R2_CONB_0;
  wire tie_lo_T3Y2__R2_CONB_0;
  wire tie_lo_T3Y30__R2_CONB_0;
  wire tie_lo_T3Y31__R2_CONB_0;
  wire tie_lo_T3Y32__R2_CONB_0;
  wire tie_lo_T3Y33__R2_CONB_0;
  wire tie_lo_T3Y34__R2_CONB_0;
  wire tie_lo_T3Y35__R2_CONB_0;
  wire tie_lo_T3Y36__R2_CONB_0;
  wire tie_lo_T3Y37__R2_CONB_0;
  wire tie_lo_T3Y38__R2_CONB_0;
  wire tie_lo_T3Y39__R2_CONB_0;
  wire tie_lo_T3Y3__R2_CONB_0;
  wire tie_lo_T3Y40__R2_CONB_0;
  wire tie_lo_T3Y41__R2_CONB_0;
  wire tie_lo_T3Y42__R2_CONB_0;
  wire tie_lo_T3Y43__R2_CONB_0;
  wire tie_lo_T3Y44__R2_CONB_0;
  wire tie_lo_T3Y45__R2_CONB_0;
  wire tie_lo_T3Y46__R2_CONB_0;
  wire tie_lo_T3Y47__R2_CONB_0;
  wire tie_lo_T3Y48__R2_CONB_0;
  wire tie_lo_T3Y49__R2_CONB_0;
  wire tie_lo_T3Y4__R2_CONB_0;
  wire tie_lo_T3Y50__R2_CONB_0;
  wire tie_lo_T3Y51__R2_CONB_0;
  wire tie_lo_T3Y52__R2_CONB_0;
  wire tie_lo_T3Y53__R2_CONB_0;
  wire tie_lo_T3Y54__R2_CONB_0;
  wire tie_lo_T3Y55__R2_CONB_0;
  wire tie_lo_T3Y56__R2_CONB_0;
  wire tie_lo_T3Y57__R2_CONB_0;
  wire tie_lo_T3Y58__R2_CONB_0;
  wire tie_lo_T3Y59__R2_CONB_0;
  wire tie_lo_T3Y5__R2_CONB_0;
  wire tie_lo_T3Y60__R2_CONB_0;
  wire tie_lo_T3Y61__R2_CONB_0;
  wire tie_lo_T3Y62__R2_CONB_0;
  wire tie_lo_T3Y63__R2_CONB_0;
  wire tie_lo_T3Y64__R2_CONB_0;
  wire tie_lo_T3Y65__R2_CONB_0;
  wire tie_lo_T3Y66__R2_CONB_0;
  wire tie_lo_T3Y67__R2_CONB_0;
  wire tie_lo_T3Y68__R2_CONB_0;
  wire tie_lo_T3Y69__R2_CONB_0;
  wire tie_lo_T3Y6__R2_CONB_0;
  wire tie_lo_T3Y70__R2_CONB_0;
  wire tie_lo_T3Y71__R2_CONB_0;
  wire tie_lo_T3Y72__R2_CONB_0;
  wire tie_lo_T3Y73__R2_CONB_0;
  wire tie_lo_T3Y74__R2_CONB_0;
  wire tie_lo_T3Y75__R2_CONB_0;
  wire tie_lo_T3Y76__R2_CONB_0;
  wire tie_lo_T3Y77__R2_CONB_0;
  wire tie_lo_T3Y78__R2_CONB_0;
  wire tie_lo_T3Y79__R2_CONB_0;
  wire tie_lo_T3Y7__R2_CONB_0;
  wire tie_lo_T3Y80__R2_CONB_0;
  wire tie_lo_T3Y81__R2_CONB_0;
  wire tie_lo_T3Y82__R2_CONB_0;
  wire tie_lo_T3Y83__R2_CONB_0;
  wire tie_lo_T3Y84__R2_CONB_0;
  wire tie_lo_T3Y85__R2_CONB_0;
  wire tie_lo_T3Y86__R2_CONB_0;
  wire tie_lo_T3Y87__R2_CONB_0;
  wire tie_lo_T3Y88__R2_CONB_0;
  wire tie_lo_T3Y89__R2_CONB_0;
  wire tie_lo_T3Y8__R2_CONB_0;
  wire tie_lo_T3Y9__R2_CONB_0;
  wire tie_lo_T4Y0__R2_CONB_0;
  wire tie_lo_T4Y10__R2_CONB_0;
  wire tie_lo_T4Y11__R2_CONB_0;
  wire tie_lo_T4Y12__R2_CONB_0;
  wire tie_lo_T4Y13__R2_CONB_0;
  wire tie_lo_T4Y14__R2_CONB_0;
  wire tie_lo_T4Y15__R2_CONB_0;
  wire tie_lo_T4Y16__R2_CONB_0;
  wire tie_lo_T4Y17__R2_CONB_0;
  wire tie_lo_T4Y18__R2_CONB_0;
  wire tie_lo_T4Y19__R2_CONB_0;
  wire tie_lo_T4Y1__R2_CONB_0;
  wire tie_lo_T4Y20__R2_CONB_0;
  wire tie_lo_T4Y21__R2_CONB_0;
  wire tie_lo_T4Y22__R2_CONB_0;
  wire tie_lo_T4Y23__R2_CONB_0;
  wire tie_lo_T4Y24__R2_CONB_0;
  wire tie_lo_T4Y25__R2_CONB_0;
  wire tie_lo_T4Y26__R2_CONB_0;
  wire tie_lo_T4Y27__R2_CONB_0;
  wire tie_lo_T4Y28__R2_CONB_0;
  wire tie_lo_T4Y29__R2_CONB_0;
  wire tie_lo_T4Y2__R2_CONB_0;
  wire tie_lo_T4Y30__R2_CONB_0;
  wire tie_lo_T4Y31__R2_CONB_0;
  wire tie_lo_T4Y32__R2_CONB_0;
  wire tie_lo_T4Y33__R2_CONB_0;
  wire tie_lo_T4Y34__R2_CONB_0;
  wire tie_lo_T4Y35__R2_CONB_0;
  wire tie_lo_T4Y36__R2_CONB_0;
  wire tie_lo_T4Y37__R2_CONB_0;
  wire tie_lo_T4Y38__R2_CONB_0;
  wire tie_lo_T4Y39__R2_CONB_0;
  wire tie_lo_T4Y3__R2_CONB_0;
  wire tie_lo_T4Y40__R2_CONB_0;
  wire tie_lo_T4Y41__R2_CONB_0;
  wire tie_lo_T4Y42__R2_CONB_0;
  wire tie_lo_T4Y43__R2_CONB_0;
  wire tie_lo_T4Y44__R2_CONB_0;
  wire tie_lo_T4Y45__R2_CONB_0;
  wire tie_lo_T4Y46__R2_CONB_0;
  wire tie_lo_T4Y47__R2_CONB_0;
  wire tie_lo_T4Y48__R2_CONB_0;
  wire tie_lo_T4Y49__R2_CONB_0;
  wire tie_lo_T4Y4__R2_CONB_0;
  wire tie_lo_T4Y50__R2_CONB_0;
  wire tie_lo_T4Y51__R2_CONB_0;
  wire tie_lo_T4Y52__R2_CONB_0;
  wire tie_lo_T4Y53__R2_CONB_0;
  wire tie_lo_T4Y54__R2_CONB_0;
  wire tie_lo_T4Y55__R2_CONB_0;
  wire tie_lo_T4Y56__R2_CONB_0;
  wire tie_lo_T4Y57__R2_CONB_0;
  wire tie_lo_T4Y58__R2_CONB_0;
  wire tie_lo_T4Y59__R2_CONB_0;
  wire tie_lo_T4Y5__R2_CONB_0;
  wire tie_lo_T4Y60__R2_CONB_0;
  wire tie_lo_T4Y61__R2_CONB_0;
  wire tie_lo_T4Y62__R2_CONB_0;
  wire tie_lo_T4Y63__R2_CONB_0;
  wire tie_lo_T4Y64__R2_CONB_0;
  wire tie_lo_T4Y65__R2_CONB_0;
  wire tie_lo_T4Y66__R2_CONB_0;
  wire tie_lo_T4Y67__R2_CONB_0;
  wire tie_lo_T4Y68__R2_CONB_0;
  wire tie_lo_T4Y69__R2_CONB_0;
  wire tie_lo_T4Y6__R2_CONB_0;
  wire tie_lo_T4Y70__R2_CONB_0;
  wire tie_lo_T4Y71__R2_CONB_0;
  wire tie_lo_T4Y72__R2_CONB_0;
  wire tie_lo_T4Y73__R2_CONB_0;
  wire tie_lo_T4Y74__R2_CONB_0;
  wire tie_lo_T4Y75__R2_CONB_0;
  wire tie_lo_T4Y76__R2_CONB_0;
  wire tie_lo_T4Y77__R2_CONB_0;
  wire tie_lo_T4Y78__R2_CONB_0;
  wire tie_lo_T4Y79__R2_CONB_0;
  wire tie_lo_T4Y7__R2_CONB_0;
  wire tie_lo_T4Y80__R2_CONB_0;
  wire tie_lo_T4Y81__R2_CONB_0;
  wire tie_lo_T4Y82__R2_CONB_0;
  wire tie_lo_T4Y83__R2_CONB_0;
  wire tie_lo_T4Y84__R2_CONB_0;
  wire tie_lo_T4Y85__R2_CONB_0;
  wire tie_lo_T4Y86__R2_CONB_0;
  wire tie_lo_T4Y87__R2_CONB_0;
  wire tie_lo_T4Y88__R2_CONB_0;
  wire tie_lo_T4Y89__R2_CONB_0;
  wire tie_lo_T4Y8__R2_CONB_0;
  wire tie_lo_T4Y9__R2_CONB_0;
  wire tie_lo_T5Y0__R2_CONB_0;
  wire tie_lo_T5Y10__R2_CONB_0;
  wire tie_lo_T5Y11__R2_CONB_0;
  wire tie_lo_T5Y12__R2_CONB_0;
  wire tie_lo_T5Y13__R2_CONB_0;
  wire tie_lo_T5Y14__R2_CONB_0;
  wire tie_lo_T5Y15__R2_CONB_0;
  wire tie_lo_T5Y16__R2_CONB_0;
  wire tie_lo_T5Y17__R2_CONB_0;
  wire tie_lo_T5Y18__R2_CONB_0;
  wire tie_lo_T5Y19__R2_CONB_0;
  wire tie_lo_T5Y1__R2_CONB_0;
  wire tie_lo_T5Y20__R2_CONB_0;
  wire tie_lo_T5Y21__R2_CONB_0;
  wire tie_lo_T5Y22__R2_CONB_0;
  wire tie_lo_T5Y23__R2_CONB_0;
  wire tie_lo_T5Y24__R2_CONB_0;
  wire tie_lo_T5Y25__R2_CONB_0;
  wire tie_lo_T5Y26__R2_CONB_0;
  wire tie_lo_T5Y27__R2_CONB_0;
  wire tie_lo_T5Y28__R2_CONB_0;
  wire tie_lo_T5Y29__R2_CONB_0;
  wire tie_lo_T5Y2__R2_CONB_0;
  wire tie_lo_T5Y30__R2_CONB_0;
  wire tie_lo_T5Y31__R2_CONB_0;
  wire tie_lo_T5Y32__R2_CONB_0;
  wire tie_lo_T5Y33__R2_CONB_0;
  wire tie_lo_T5Y34__R2_CONB_0;
  wire tie_lo_T5Y35__R2_CONB_0;
  wire tie_lo_T5Y36__R2_CONB_0;
  wire tie_lo_T5Y37__R2_CONB_0;
  wire tie_lo_T5Y38__R2_CONB_0;
  wire tie_lo_T5Y39__R2_CONB_0;
  wire tie_lo_T5Y3__R2_CONB_0;
  wire tie_lo_T5Y40__R2_CONB_0;
  wire tie_lo_T5Y41__R2_CONB_0;
  wire tie_lo_T5Y42__R2_CONB_0;
  wire tie_lo_T5Y43__R2_CONB_0;
  wire tie_lo_T5Y44__R2_CONB_0;
  wire tie_lo_T5Y45__R2_CONB_0;
  wire tie_lo_T5Y46__R2_CONB_0;
  wire tie_lo_T5Y47__R2_CONB_0;
  wire tie_lo_T5Y48__R2_CONB_0;
  wire tie_lo_T5Y49__R2_CONB_0;
  wire tie_lo_T5Y4__R2_CONB_0;
  wire tie_lo_T5Y50__R2_CONB_0;
  wire tie_lo_T5Y51__R2_CONB_0;
  wire tie_lo_T5Y52__R2_CONB_0;
  wire tie_lo_T5Y53__R2_CONB_0;
  wire tie_lo_T5Y54__R2_CONB_0;
  wire tie_lo_T5Y55__R2_CONB_0;
  wire tie_lo_T5Y56__R2_CONB_0;
  wire tie_lo_T5Y57__R2_CONB_0;
  wire tie_lo_T5Y58__R2_CONB_0;
  wire tie_lo_T5Y59__R2_CONB_0;
  wire tie_lo_T5Y5__R2_CONB_0;
  wire tie_lo_T5Y60__R2_CONB_0;
  wire tie_lo_T5Y61__R2_CONB_0;
  wire tie_lo_T5Y62__R2_CONB_0;
  wire tie_lo_T5Y63__R2_CONB_0;
  wire tie_lo_T5Y64__R2_CONB_0;
  wire tie_lo_T5Y65__R2_CONB_0;
  wire tie_lo_T5Y66__R2_CONB_0;
  wire tie_lo_T5Y67__R2_CONB_0;
  wire tie_lo_T5Y68__R2_CONB_0;
  wire tie_lo_T5Y69__R2_CONB_0;
  wire tie_lo_T5Y6__R2_CONB_0;
  wire tie_lo_T5Y70__R2_CONB_0;
  wire tie_lo_T5Y71__R2_CONB_0;
  wire tie_lo_T5Y72__R2_CONB_0;
  wire tie_lo_T5Y73__R2_CONB_0;
  wire tie_lo_T5Y74__R2_CONB_0;
  wire tie_lo_T5Y75__R2_CONB_0;
  wire tie_lo_T5Y76__R2_CONB_0;
  wire tie_lo_T5Y77__R2_CONB_0;
  wire tie_lo_T5Y78__R2_CONB_0;
  wire tie_lo_T5Y79__R2_CONB_0;
  wire tie_lo_T5Y7__R2_CONB_0;
  wire tie_lo_T5Y80__R2_CONB_0;
  wire tie_lo_T5Y81__R2_CONB_0;
  wire tie_lo_T5Y82__R2_CONB_0;
  wire tie_lo_T5Y83__R2_CONB_0;
  wire tie_lo_T5Y84__R2_CONB_0;
  wire tie_lo_T5Y85__R2_CONB_0;
  wire tie_lo_T5Y86__R2_CONB_0;
  wire tie_lo_T5Y87__R2_CONB_0;
  wire tie_lo_T5Y88__R2_CONB_0;
  wire tie_lo_T5Y89__R2_CONB_0;
  wire tie_lo_T5Y8__R2_CONB_0;
  wire tie_lo_T5Y9__R2_CONB_0;
  wire tie_lo_T6Y0__R2_CONB_0;
  wire tie_lo_T6Y10__R2_CONB_0;
  wire tie_lo_T6Y11__R2_CONB_0;
  wire tie_lo_T6Y12__R2_CONB_0;
  wire tie_lo_T6Y13__R2_CONB_0;
  wire tie_lo_T6Y14__R2_CONB_0;
  wire tie_lo_T6Y15__R2_CONB_0;
  wire tie_lo_T6Y16__R2_CONB_0;
  wire tie_lo_T6Y17__R2_CONB_0;
  wire tie_lo_T6Y18__R2_CONB_0;
  wire tie_lo_T6Y19__R2_CONB_0;
  wire tie_lo_T6Y1__R2_CONB_0;
  wire tie_lo_T6Y20__R2_CONB_0;
  wire tie_lo_T6Y21__R2_CONB_0;
  wire tie_lo_T6Y22__R2_CONB_0;
  wire tie_lo_T6Y23__R2_CONB_0;
  wire tie_lo_T6Y24__R2_CONB_0;
  wire tie_lo_T6Y25__R2_CONB_0;
  wire tie_lo_T6Y26__R2_CONB_0;
  wire tie_lo_T6Y27__R2_CONB_0;
  wire tie_lo_T6Y28__R2_CONB_0;
  wire tie_lo_T6Y29__R2_CONB_0;
  wire tie_lo_T6Y2__R2_CONB_0;
  wire tie_lo_T6Y30__R2_CONB_0;
  wire tie_lo_T6Y31__R2_CONB_0;
  wire tie_lo_T6Y32__R2_CONB_0;
  wire tie_lo_T6Y33__R2_CONB_0;
  wire tie_lo_T6Y34__R2_CONB_0;
  wire tie_lo_T6Y35__R2_CONB_0;
  wire tie_lo_T6Y36__R2_CONB_0;
  wire tie_lo_T6Y37__R2_CONB_0;
  wire tie_lo_T6Y38__R2_CONB_0;
  wire tie_lo_T6Y39__R2_CONB_0;
  wire tie_lo_T6Y3__R2_CONB_0;
  wire tie_lo_T6Y40__R2_CONB_0;
  wire tie_lo_T6Y41__R2_CONB_0;
  wire tie_lo_T6Y42__R2_CONB_0;
  wire tie_lo_T6Y43__R2_CONB_0;
  wire tie_lo_T6Y44__R2_CONB_0;
  wire tie_lo_T6Y45__R2_CONB_0;
  wire tie_lo_T6Y46__R2_CONB_0;
  wire tie_lo_T6Y47__R2_CONB_0;
  wire tie_lo_T6Y48__R2_CONB_0;
  wire tie_lo_T6Y49__R2_CONB_0;
  wire tie_lo_T6Y4__R2_CONB_0;
  wire tie_lo_T6Y50__R2_CONB_0;
  wire tie_lo_T6Y51__R2_CONB_0;
  wire tie_lo_T6Y52__R2_CONB_0;
  wire tie_lo_T6Y53__R2_CONB_0;
  wire tie_lo_T6Y54__R2_CONB_0;
  wire tie_lo_T6Y55__R2_CONB_0;
  wire tie_lo_T6Y56__R2_CONB_0;
  wire tie_lo_T6Y57__R2_CONB_0;
  wire tie_lo_T6Y58__R2_CONB_0;
  wire tie_lo_T6Y59__R2_CONB_0;
  wire tie_lo_T6Y5__R2_CONB_0;
  wire tie_lo_T6Y60__R2_CONB_0;
  wire tie_lo_T6Y61__R2_CONB_0;
  wire tie_lo_T6Y62__R2_CONB_0;
  wire tie_lo_T6Y63__R2_CONB_0;
  wire tie_lo_T6Y64__R2_CONB_0;
  wire tie_lo_T6Y65__R2_CONB_0;
  wire tie_lo_T6Y66__R2_CONB_0;
  wire tie_lo_T6Y67__R2_CONB_0;
  wire tie_lo_T6Y68__R2_CONB_0;
  wire tie_lo_T6Y69__R2_CONB_0;
  wire tie_lo_T6Y6__R2_CONB_0;
  wire tie_lo_T6Y70__R2_CONB_0;
  wire tie_lo_T6Y71__R2_CONB_0;
  wire tie_lo_T6Y72__R2_CONB_0;
  wire tie_lo_T6Y73__R2_CONB_0;
  wire tie_lo_T6Y74__R2_CONB_0;
  wire tie_lo_T6Y75__R2_CONB_0;
  wire tie_lo_T6Y76__R2_CONB_0;
  wire tie_lo_T6Y77__R2_CONB_0;
  wire tie_lo_T6Y78__R2_CONB_0;
  wire tie_lo_T6Y79__R2_CONB_0;
  wire tie_lo_T6Y7__R2_CONB_0;
  wire tie_lo_T6Y80__R2_CONB_0;
  wire tie_lo_T6Y81__R2_CONB_0;
  wire tie_lo_T6Y82__R2_CONB_0;
  wire tie_lo_T6Y83__R2_CONB_0;
  wire tie_lo_T6Y84__R2_CONB_0;
  wire tie_lo_T6Y85__R2_CONB_0;
  wire tie_lo_T6Y86__R2_CONB_0;
  wire tie_lo_T6Y87__R2_CONB_0;
  wire tie_lo_T6Y88__R2_CONB_0;
  wire tie_lo_T6Y89__R2_CONB_0;
  wire tie_lo_T6Y8__R2_CONB_0;
  wire tie_lo_T6Y9__R2_CONB_0;
  wire tie_lo_T7Y0__R2_CONB_0;
  wire tie_lo_T7Y10__R2_CONB_0;
  wire tie_lo_T7Y11__R2_CONB_0;
  wire tie_lo_T7Y12__R2_CONB_0;
  wire tie_lo_T7Y13__R2_CONB_0;
  wire tie_lo_T7Y14__R2_CONB_0;
  wire tie_lo_T7Y15__R2_CONB_0;
  wire tie_lo_T7Y16__R2_CONB_0;
  wire tie_lo_T7Y17__R2_CONB_0;
  wire tie_lo_T7Y18__R2_CONB_0;
  wire tie_lo_T7Y19__R2_CONB_0;
  wire tie_lo_T7Y1__R2_CONB_0;
  wire tie_lo_T7Y20__R2_CONB_0;
  wire tie_lo_T7Y21__R2_CONB_0;
  wire tie_lo_T7Y22__R2_CONB_0;
  wire tie_lo_T7Y23__R2_CONB_0;
  wire tie_lo_T7Y24__R2_CONB_0;
  wire tie_lo_T7Y25__R2_CONB_0;
  wire tie_lo_T7Y26__R2_CONB_0;
  wire tie_lo_T7Y27__R2_CONB_0;
  wire tie_lo_T7Y28__R2_CONB_0;
  wire tie_lo_T7Y29__R2_CONB_0;
  wire tie_lo_T7Y2__R2_CONB_0;
  wire tie_lo_T7Y30__R2_CONB_0;
  wire tie_lo_T7Y31__R2_CONB_0;
  wire tie_lo_T7Y32__R2_CONB_0;
  wire tie_lo_T7Y33__R2_CONB_0;
  wire tie_lo_T7Y34__R2_CONB_0;
  wire tie_lo_T7Y35__R2_CONB_0;
  wire tie_lo_T7Y36__R2_CONB_0;
  wire tie_lo_T7Y37__R2_CONB_0;
  wire tie_lo_T7Y38__R2_CONB_0;
  wire tie_lo_T7Y39__R2_CONB_0;
  wire tie_lo_T7Y3__R2_CONB_0;
  wire tie_lo_T7Y40__R2_CONB_0;
  wire tie_lo_T7Y41__R2_CONB_0;
  wire tie_lo_T7Y42__R2_CONB_0;
  wire tie_lo_T7Y43__R2_CONB_0;
  wire tie_lo_T7Y44__R2_CONB_0;
  wire tie_lo_T7Y45__R2_CONB_0;
  wire tie_lo_T7Y46__R2_CONB_0;
  wire tie_lo_T7Y47__R2_CONB_0;
  wire tie_lo_T7Y48__R2_CONB_0;
  wire tie_lo_T7Y49__R2_CONB_0;
  wire tie_lo_T7Y4__R2_CONB_0;
  wire tie_lo_T7Y50__R2_CONB_0;
  wire tie_lo_T7Y51__R2_CONB_0;
  wire tie_lo_T7Y52__R2_CONB_0;
  wire tie_lo_T7Y53__R2_CONB_0;
  wire tie_lo_T7Y54__R2_CONB_0;
  wire tie_lo_T7Y55__R2_CONB_0;
  wire tie_lo_T7Y56__R2_CONB_0;
  wire tie_lo_T7Y57__R2_CONB_0;
  wire tie_lo_T7Y58__R2_CONB_0;
  wire tie_lo_T7Y59__R2_CONB_0;
  wire tie_lo_T7Y5__R2_CONB_0;
  wire tie_lo_T7Y60__R2_CONB_0;
  wire tie_lo_T7Y61__R2_CONB_0;
  wire tie_lo_T7Y62__R2_CONB_0;
  wire tie_lo_T7Y63__R2_CONB_0;
  wire tie_lo_T7Y64__R2_CONB_0;
  wire tie_lo_T7Y65__R2_CONB_0;
  wire tie_lo_T7Y66__R2_CONB_0;
  wire tie_lo_T7Y67__R2_CONB_0;
  wire tie_lo_T7Y68__R2_CONB_0;
  wire tie_lo_T7Y69__R2_CONB_0;
  wire tie_lo_T7Y6__R2_CONB_0;
  wire tie_lo_T7Y70__R2_CONB_0;
  wire tie_lo_T7Y71__R2_CONB_0;
  wire tie_lo_T7Y72__R2_CONB_0;
  wire tie_lo_T7Y73__R2_CONB_0;
  wire tie_lo_T7Y74__R2_CONB_0;
  wire tie_lo_T7Y75__R2_CONB_0;
  wire tie_lo_T7Y76__R2_CONB_0;
  wire tie_lo_T7Y77__R2_CONB_0;
  wire tie_lo_T7Y78__R2_CONB_0;
  wire tie_lo_T7Y79__R2_CONB_0;
  wire tie_lo_T7Y7__R2_CONB_0;
  wire tie_lo_T7Y80__R2_CONB_0;
  wire tie_lo_T7Y81__R2_CONB_0;
  wire tie_lo_T7Y82__R2_CONB_0;
  wire tie_lo_T7Y83__R2_CONB_0;
  wire tie_lo_T7Y84__R2_CONB_0;
  wire tie_lo_T7Y85__R2_CONB_0;
  wire tie_lo_T7Y86__R2_CONB_0;
  wire tie_lo_T7Y87__R2_CONB_0;
  wire tie_lo_T7Y88__R2_CONB_0;
  wire tie_lo_T7Y89__R2_CONB_0;
  wire tie_lo_T7Y8__R2_CONB_0;
  wire tie_lo_T7Y9__R2_CONB_0;
  wire tie_lo_T8Y0__R2_CONB_0;
  wire tie_lo_T8Y10__R2_CONB_0;
  wire tie_lo_T8Y11__R2_CONB_0;
  wire tie_lo_T8Y12__R2_CONB_0;
  wire tie_lo_T8Y13__R2_CONB_0;
  wire tie_lo_T8Y14__R2_CONB_0;
  wire tie_lo_T8Y15__R2_CONB_0;
  wire tie_lo_T8Y16__R2_CONB_0;
  wire tie_lo_T8Y17__R2_CONB_0;
  wire tie_lo_T8Y18__R2_CONB_0;
  wire tie_lo_T8Y19__R2_CONB_0;
  wire tie_lo_T8Y1__R2_CONB_0;
  wire tie_lo_T8Y20__R2_CONB_0;
  wire tie_lo_T8Y21__R2_CONB_0;
  wire tie_lo_T8Y22__R2_CONB_0;
  wire tie_lo_T8Y23__R2_CONB_0;
  wire tie_lo_T8Y24__R2_CONB_0;
  wire tie_lo_T8Y25__R2_CONB_0;
  wire tie_lo_T8Y26__R2_CONB_0;
  wire tie_lo_T8Y27__R2_CONB_0;
  wire tie_lo_T8Y28__R2_CONB_0;
  wire tie_lo_T8Y29__R2_CONB_0;
  wire tie_lo_T8Y2__R2_CONB_0;
  wire tie_lo_T8Y30__R2_CONB_0;
  wire tie_lo_T8Y31__R2_CONB_0;
  wire tie_lo_T8Y32__R2_CONB_0;
  wire tie_lo_T8Y33__R2_CONB_0;
  wire tie_lo_T8Y34__R2_CONB_0;
  wire tie_lo_T8Y35__R2_CONB_0;
  wire tie_lo_T8Y36__R2_CONB_0;
  wire tie_lo_T8Y37__R2_CONB_0;
  wire tie_lo_T8Y38__R2_CONB_0;
  wire tie_lo_T8Y39__R2_CONB_0;
  wire tie_lo_T8Y3__R2_CONB_0;
  wire tie_lo_T8Y40__R2_CONB_0;
  wire tie_lo_T8Y41__R2_CONB_0;
  wire tie_lo_T8Y42__R2_CONB_0;
  wire tie_lo_T8Y43__R2_CONB_0;
  wire tie_lo_T8Y44__R2_CONB_0;
  wire tie_lo_T8Y45__R2_CONB_0;
  wire tie_lo_T8Y46__R2_CONB_0;
  wire tie_lo_T8Y47__R2_CONB_0;
  wire tie_lo_T8Y48__R2_CONB_0;
  wire tie_lo_T8Y49__R2_CONB_0;
  wire tie_lo_T8Y4__R2_CONB_0;
  wire tie_lo_T8Y50__R2_CONB_0;
  wire tie_lo_T8Y51__R2_CONB_0;
  wire tie_lo_T8Y52__R2_CONB_0;
  wire tie_lo_T8Y53__R2_CONB_0;
  wire tie_lo_T8Y54__R2_CONB_0;
  wire tie_lo_T8Y55__R2_CONB_0;
  wire tie_lo_T8Y56__R2_CONB_0;
  wire tie_lo_T8Y57__R2_CONB_0;
  wire tie_lo_T8Y58__R2_CONB_0;
  wire tie_lo_T8Y59__R2_CONB_0;
  wire tie_lo_T8Y5__R2_CONB_0;
  wire tie_lo_T8Y60__R2_CONB_0;
  wire tie_lo_T8Y61__R2_CONB_0;
  wire tie_lo_T8Y62__R2_CONB_0;
  wire tie_lo_T8Y63__R2_CONB_0;
  wire tie_lo_T8Y64__R2_CONB_0;
  wire tie_lo_T8Y65__R2_CONB_0;
  wire tie_lo_T8Y66__R2_CONB_0;
  wire tie_lo_T8Y67__R2_CONB_0;
  wire tie_lo_T8Y68__R2_CONB_0;
  wire tie_lo_T8Y69__R2_CONB_0;
  wire tie_lo_T8Y6__R2_CONB_0;
  wire tie_lo_T8Y70__R2_CONB_0;
  wire tie_lo_T8Y71__R2_CONB_0;
  wire tie_lo_T8Y72__R2_CONB_0;
  wire tie_lo_T8Y73__R2_CONB_0;
  wire tie_lo_T8Y74__R2_CONB_0;
  wire tie_lo_T8Y75__R2_CONB_0;
  wire tie_lo_T8Y76__R2_CONB_0;
  wire tie_lo_T8Y77__R2_CONB_0;
  wire tie_lo_T8Y78__R2_CONB_0;
  wire tie_lo_T8Y79__R2_CONB_0;
  wire tie_lo_T8Y7__R2_CONB_0;
  wire tie_lo_T8Y80__R2_CONB_0;
  wire tie_lo_T8Y81__R2_CONB_0;
  wire tie_lo_T8Y82__R2_CONB_0;
  wire tie_lo_T8Y83__R2_CONB_0;
  wire tie_lo_T8Y84__R2_CONB_0;
  wire tie_lo_T8Y85__R2_CONB_0;
  wire tie_lo_T8Y86__R2_CONB_0;
  wire tie_lo_T8Y87__R2_CONB_0;
  wire tie_lo_T8Y88__R2_CONB_0;
  wire tie_lo_T8Y89__R2_CONB_0;
  wire tie_lo_T8Y8__R2_CONB_0;
  wire tie_lo_T8Y9__R2_CONB_0;
  wire tie_lo_T9Y0__R2_CONB_0;
  wire tie_lo_T9Y10__R2_CONB_0;
  wire tie_lo_T9Y11__R2_CONB_0;
  wire tie_lo_T9Y12__R2_CONB_0;
  wire tie_lo_T9Y13__R2_CONB_0;
  wire tie_lo_T9Y14__R2_CONB_0;
  wire tie_lo_T9Y15__R2_CONB_0;
  wire tie_lo_T9Y16__R2_CONB_0;
  wire tie_lo_T9Y17__R2_CONB_0;
  wire tie_lo_T9Y18__R2_CONB_0;
  wire tie_lo_T9Y19__R2_CONB_0;
  wire tie_lo_T9Y1__R2_CONB_0;
  wire tie_lo_T9Y20__R2_CONB_0;
  wire tie_lo_T9Y21__R2_CONB_0;
  wire tie_lo_T9Y22__R2_CONB_0;
  wire tie_lo_T9Y23__R2_CONB_0;
  wire tie_lo_T9Y24__R2_CONB_0;
  wire tie_lo_T9Y25__R2_CONB_0;
  wire tie_lo_T9Y26__R2_CONB_0;
  wire tie_lo_T9Y27__R2_CONB_0;
  wire tie_lo_T9Y28__R2_CONB_0;
  wire tie_lo_T9Y29__R2_CONB_0;
  wire tie_lo_T9Y2__R2_CONB_0;
  wire tie_lo_T9Y30__R2_CONB_0;
  wire tie_lo_T9Y31__R2_CONB_0;
  wire tie_lo_T9Y32__R2_CONB_0;
  wire tie_lo_T9Y33__R2_CONB_0;
  wire tie_lo_T9Y34__R2_CONB_0;
  wire tie_lo_T9Y35__R2_CONB_0;
  wire tie_lo_T9Y36__R2_CONB_0;
  wire tie_lo_T9Y37__R2_CONB_0;
  wire tie_lo_T9Y38__R2_CONB_0;
  wire tie_lo_T9Y39__R2_CONB_0;
  wire tie_lo_T9Y3__R2_CONB_0;
  wire tie_lo_T9Y40__R2_CONB_0;
  wire tie_lo_T9Y41__R2_CONB_0;
  wire tie_lo_T9Y42__R2_CONB_0;
  wire tie_lo_T9Y43__R2_CONB_0;
  wire tie_lo_T9Y44__R2_CONB_0;
  wire tie_lo_T9Y45__R2_CONB_0;
  wire tie_lo_T9Y46__R2_CONB_0;
  wire tie_lo_T9Y47__R2_CONB_0;
  wire tie_lo_T9Y48__R2_CONB_0;
  wire tie_lo_T9Y49__R2_CONB_0;
  wire tie_lo_T9Y4__R2_CONB_0;
  wire tie_lo_T9Y50__R2_CONB_0;
  wire tie_lo_T9Y51__R2_CONB_0;
  wire tie_lo_T9Y52__R2_CONB_0;
  wire tie_lo_T9Y53__R2_CONB_0;
  wire tie_lo_T9Y54__R2_CONB_0;
  wire tie_lo_T9Y55__R2_CONB_0;
  wire tie_lo_T9Y56__R2_CONB_0;
  wire tie_lo_T9Y57__R2_CONB_0;
  wire tie_lo_T9Y58__R2_CONB_0;
  wire tie_lo_T9Y59__R2_CONB_0;
  wire tie_lo_T9Y5__R2_CONB_0;
  wire tie_lo_T9Y60__R2_CONB_0;
  wire tie_lo_T9Y61__R2_CONB_0;
  wire tie_lo_T9Y62__R2_CONB_0;
  wire tie_lo_T9Y63__R2_CONB_0;
  wire tie_lo_T9Y64__R2_CONB_0;
  wire tie_lo_T9Y65__R2_CONB_0;
  wire tie_lo_T9Y66__R2_CONB_0;
  wire tie_lo_T9Y67__R2_CONB_0;
  wire tie_lo_T9Y68__R2_CONB_0;
  wire tie_lo_T9Y69__R2_CONB_0;
  wire tie_lo_T9Y6__R2_CONB_0;
  wire tie_lo_T9Y70__R2_CONB_0;
  wire tie_lo_T9Y71__R2_CONB_0;
  wire tie_lo_T9Y72__R2_CONB_0;
  wire tie_lo_T9Y73__R2_CONB_0;
  wire tie_lo_T9Y74__R2_CONB_0;
  wire tie_lo_T9Y75__R2_CONB_0;
  wire tie_lo_T9Y76__R2_CONB_0;
  wire tie_lo_T9Y77__R2_CONB_0;
  wire tie_lo_T9Y78__R2_CONB_0;
  wire tie_lo_T9Y79__R2_CONB_0;
  wire tie_lo_T9Y7__R2_CONB_0;
  wire tie_lo_T9Y80__R2_CONB_0;
  wire tie_lo_T9Y81__R2_CONB_0;
  wire tie_lo_T9Y82__R2_CONB_0;
  wire tie_lo_T9Y83__R2_CONB_0;
  wire tie_lo_T9Y84__R2_CONB_0;
  wire tie_lo_T9Y85__R2_CONB_0;
  wire tie_lo_T9Y86__R2_CONB_0;
  wire tie_lo_T9Y87__R2_CONB_0;
  wire tie_lo_T9Y88__R2_CONB_0;
  wire tie_lo_T9Y89__R2_CONB_0;
  wire tie_lo_T9Y8__R2_CONB_0;
  wire tie_lo_T9Y9__R2_CONB_0;

  // Cell instantiations
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10000 (.A([124]), .B([125]), .X([126]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10001 (.A([127]), .B([126]), .X([128]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10002 (.A([128]), .Y([129]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10003 (.A([130]), .B([129]), .Y([131]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10004 (.A([132]), .B([131]), .Y([133]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10005 (.A([133]), .Y([134]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10006 (.A([132]), .B([131]), .X([135]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10007 (.A([133]), .B([135]), .Y([136]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10008 (.A([39]), .B([136]), .Y([137]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10009 (.A([39]), .B([138]), .X([139]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10010 (.A([137]), .B([139]), .Y([140]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10011 (.A([140]), .Y([141]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10012 (.A([142]), .B([143]), .Y([144]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10013 (.A([145]), .B([146]), .Y([147]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10014 (.A([145]), .B([148]), .Y([149]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10015 (.A([150]), .B([149]), .Y([151]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10016 (.A([152]), .B([153]), .Y([154]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10017 (.A([147]), .B([154]), .Y([155]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10018 (.A([151]), .B([155]), .X([156]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10019 (.A([156]), .Y([157]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10020 (.A([144]), .B([157]), .Y([158]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10021 (.A([134]), .B([158]), .Y([159]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10022 (.A([159]), .Y([160]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10023 (.A([134]), .B([158]), .X([161]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10024 (.A([159]), .B([161]), .Y([162]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10025 (.A([39]), .B([162]), .Y([163]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10026 (.A([39]), .B([142]), .X([164]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10027 (.A([163]), .B([164]), .Y([165]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10028 (.A([165]), .Y([166]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10029 (.A([167]), .B([143]), .Y([168]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10030 (.A([169]), .B([146]), .Y([170]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10031 (.A([171]), .B([172]), .X([173]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10032 (.A([150]), .B([173]), .Y([174]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10033 (.A([175]), .B([153]), .Y([176]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10034 (.A([170]), .B([176]), .Y([177]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10035 (.A([174]), .B([177]), .X([178]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10036 (.A([178]), .Y([179]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10037 (.A([168]), .B([179]), .Y([180]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10038 (.A([160]), .B([180]), .Y([181]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10039 (.A([181]), .Y([182]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10040 (.A([160]), .B([180]), .X([183]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10041 (.A([181]), .B([183]), .Y([184]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10042 (.A([39]), .B([184]), .Y([185]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10043 (.A([39]), .B([167]), .X([186]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10044 (.A([185]), .B([186]), .Y([187]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10045 (.A([187]), .Y([188]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10046 (.A([189]), .B([143]), .Y([190]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10047 (.A([191]), .B([146]), .Y([192]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10048 (.A([191]), .B([148]), .Y([193]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10049 (.A([194]), .B([153]), .Y([195]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10050 (.A([193]), .B([195]), .Y([196]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10051 (.A([196]), .Y([197]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10052 (.A([192]), .B([197]), .Y([198]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10053 (.A([199]), .B([198]), .X([200]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10054 (.A([200]), .Y([201]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10055 (.A([190]), .B([201]), .Y([202]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10056 (.A([182]), .B([202]), .Y([203]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10057 (.A([203]), .Y([204]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10058 (.A([182]), .B([202]), .X([205]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10059 (.A([203]), .B([205]), .Y([206]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10060 (.A([39]), .B([189]), .X([207]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10061 (.A([39]), .B([206]), .Y([208]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10062 (.A([207]), .B([208]), .Y([209]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10063 (.A([209]), .Y([210]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10064 (.A([211]), .B([143]), .Y([212]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10065 (.A([213]), .B([146]), .Y([214]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10066 (.A([215]), .B([172]), .X([216]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10067 (.A([150]), .B([216]), .Y([217]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10068 (.A([218]), .B([153]), .Y([219]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10069 (.A([214]), .B([219]), .Y([220]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10070 (.A([217]), .B([220]), .X([221]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10071 (.A([221]), .Y([222]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10072 (.A([212]), .B([222]), .Y([223]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10073 (.A([204]), .B([223]), .Y([224]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10074 (.A([224]), .Y([225]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10075 (.A([204]), .B([223]), .X([226]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10076 (.A([224]), .B([226]), .Y([227]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10077 (.A([39]), .B([227]), .Y([228]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10078 (.A([39]), .B([211]), .X([229]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10079 (.A([228]), .B([229]), .Y([230]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10080 (.A([230]), .Y([231]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10081 (.A([232]), .B([143]), .Y([233]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10082 (.A([234]), .B([146]), .Y([235]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10083 (.A([236]), .B([172]), .X([237]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10084 (.A([150]), .B([237]), .Y([238]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10085 (.A([239]), .B([153]), .Y([240]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10086 (.A([235]), .B([240]), .Y([241]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10087 (.A([238]), .B([241]), .X([242]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10088 (.A([242]), .Y([243]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10089 (.A([233]), .B([243]), .Y([244]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10090 (.A([225]), .B([244]), .Y([245]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10091 (.A([245]), .Y([246]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10092 (.A([225]), .B([244]), .X([247]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10093 (.A([245]), .B([247]), .Y([248]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10094 (.A([39]), .B([232]), .X([249]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10095 (.A([39]), .B([248]), .Y([250]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10096 (.A([249]), .B([250]), .Y([251]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10097 (.A([251]), .Y([252]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10098 (.A([253]), .B([254]), .Y([255]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10099 (.A([256]), .B([146]), .Y([257]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10100 (.A([258]), .B([153]), .Y([259]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10101 (.A([258]), .B([148]), .Y([260]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10102 (.A([150]), .B([260]), .Y([261]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10103 (.A([261]), .Y([262]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10104 (.A([263]), .B([264]), .X([265]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10105 (.A([259]), .B([262]), .Y([266]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10106 (.A([257]), .B([265]), .Y([267]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10107 (.A([266]), .B([267]), .X([268]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10108 (.A([268]), .Y([269]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10109 (.A([255]), .B([269]), .Y([270]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10110 (.A([246]), .B([270]), .Y([271]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10111 (.A([271]), .Y([272]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10112 (.A([246]), .B([270]), .X([273]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10113 (.A([271]), .B([273]), .Y([274]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10114 (.A([39]), .B([274]), .Y([275]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10115 (.A([39]), .B([253]), .X([276]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10116 (.A([275]), .B([276]), .Y([277]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10117 (.A([277]), .Y([278]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10118 (.A([279]), .B([254]), .Y([280]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10119 (.A([281]), .B([146]), .Y([282]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10120 (.A([283]), .B([153]), .Y([284]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10121 (.A([283]), .B([148]), .Y([285]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10122 (.A([286]), .B([287]), .Y([288]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10123 (.A([284]), .B([285]), .Y([289]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10124 (.A([199]), .B([289]), .X([290]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10125 (.A([282]), .B([288]), .Y([291]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10126 (.A([290]), .B([291]), .X([292]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10127 (.A([292]), .Y([293]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10128 (.A([280]), .B([293]), .Y([294]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10129 (.A([272]), .B([294]), .Y([295]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10130 (.A([295]), .Y([296]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10131 (.A([272]), .B([294]), .X([297]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10132 (.A([295]), .B([297]), .Y([298]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10133 (.A([39]), .B([298]), .Y([299]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10134 (.A([39]), .B([279]), .X([300]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10135 (.A([299]), .B([300]), .Y([301]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10136 (.A([301]), .Y([302]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10137 (.A([303]), .B([254]), .Y([304]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10138 (.A([305]), .B([146]), .Y([306]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10139 (.A([307]), .B([153]), .Y([308]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10140 (.A([309]), .B([264]), .X([310]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10141 (.A([307]), .B([148]), .Y([311]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10142 (.A([311]), .Y([312]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10143 (.A([150]), .B([308]), .Y([313]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10144 (.A([312]), .B([313]), .X([314]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10145 (.A([306]), .B([310]), .Y([315]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10146 (.A([314]), .B([315]), .X([316]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10147 (.A([316]), .Y([317]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10148 (.A([304]), .B([317]), .Y([318]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10149 (.A([296]), .B([318]), .Y([319]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10150 (.A([319]), .Y([320]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10151 (.A([296]), .B([318]), .X([321]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10152 (.A([319]), .B([321]), .Y([322]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10153 (.A([39]), .B([303]), .X([323]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10154 (.A([39]), .B([322]), .Y([324]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10155 (.A([323]), .B([324]), .Y([325]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10156 (.A([325]), .Y([326]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10157 (.A([327]), .B([254]), .Y([328]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10158 (.A([329]), .B([146]), .Y([330]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10159 (.A([331]), .B([153]), .Y([332]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10160 (.A([145]), .B([287]), .Y([333]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10161 (.A([331]), .B([148]), .Y([334]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10162 (.A([333]), .B([334]), .Y([335]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10163 (.A([199]), .B([335]), .X([336]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10164 (.A([330]), .B([332]), .Y([337]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10165 (.A([336]), .B([337]), .X([338]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10166 (.A([338]), .Y([339]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10167 (.A([328]), .B([339]), .Y([340]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10168 (.A([320]), .B([340]), .Y([341]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10169 (.A([341]), .Y([342]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10170 (.A([320]), .B([340]), .X([343]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10171 (.A([341]), .B([343]), .Y([344]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10172 (.A([39]), .B([344]), .Y([345]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10173 (.A([39]), .B([327]), .X([346]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10174 (.A([345]), .B([346]), .Y([347]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10175 (.A([347]), .Y([348]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10176 (.A([349]), .B([254]), .Y([350]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10177 (.A([350]), .Y([351]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10178 (.A([352]), .B([146]), .Y([353]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10179 (.A([353]), .Y([354]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10180 (.A([355]), .B([153]), .Y([356]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10181 (.A([171]), .B([264]), .X([357]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10182 (.A([355]), .B([148]), .Y([358]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10183 (.A([358]), .Y([359]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10184 (.A([356]), .B([357]), .Y([360]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10185 (.A([359]), .B([360]), .X([361]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10186 (.A([354]), .B([361]), .X([362]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10187 (.A([199]), .B([362]), .X([363]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10188 (.A([351]), .B([363]), .X([364]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10189 (.A([342]), .B([364]), .Y([365]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10190 (.A([365]), .Y([366]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10191 (.A([342]), .B([364]), .X([367]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10192 (.A([365]), .B([367]), .Y([368]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10193 (.A([39]), .B([368]), .Y([369]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10194 (.A([39]), .B([349]), .X([370]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10195 (.A([369]), .B([370]), .Y([371]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10196 (.A([371]), .Y([372]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10197 (.A([373]), .B([254]), .Y([374]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10198 (.A([375]), .B([146]), .Y([376]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10199 (.A([376]), .Y([377]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10200 (.A([378]), .B([153]), .Y([379]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10201 (.A([378]), .B([148]), .Y([380]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10202 (.A([150]), .B([380]), .Y([381]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10203 (.A([191]), .B([287]), .Y([382]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10204 (.A([379]), .B([382]), .Y([383]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10205 (.A([381]), .B([383]), .X([384]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10206 (.A([384]), .Y([385]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10207 (.A([374]), .B([385]), .Y([386]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10208 (.A([377]), .B([386]), .X([387]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10209 (.A([366]), .B([387]), .Y([388]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10210 (.A([388]), .Y([389]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10211 (.A([366]), .B([387]), .X([390]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10212 (.A([388]), .B([390]), .Y([391]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10213 (.A([39]), .B([391]), .Y([392]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10214 (.A([39]), .B([373]), .X([393]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10215 (.A([392]), .B([393]), .Y([394]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10216 (.A([394]), .Y([395]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10217 (.A([396]), .B([254]), .Y([397]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10218 (.A([398]), .B([146]), .Y([399]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10219 (.A([400]), .B([148]), .Y([401]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10220 (.A([215]), .B([264]), .X([402]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10221 (.A([401]), .B([402]), .Y([403]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10222 (.A([199]), .B([403]), .X([404]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10223 (.A([400]), .B([153]), .Y([405]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10224 (.A([399]), .B([405]), .Y([406]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10225 (.A([404]), .B([406]), .X([407]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10226 (.A([407]), .Y([408]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10227 (.A([397]), .B([408]), .Y([409]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10228 (.A([389]), .B([409]), .Y([410]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10229 (.A([389]), .B([409]), .X([411]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10230 (.A([410]), .B([411]), .Y([412]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10231 (.A([39]), .B([412]), .Y([413]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10232 (.A([39]), .B([396]), .X([414]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10233 (.A([413]), .B([414]), .Y([415]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10234 (.A([415]), .Y([416]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10235 (.A([417]), .B([254]), .Y([418]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10236 (.A([419]), .B([146]), .Y([420]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10237 (.A([421]), .B([153]), .Y([422]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10238 (.A([236]), .B([264]), .X([423]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10239 (.A([421]), .B([148]), .Y([424]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10240 (.A([420]), .B([423]), .Y([425]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10241 (.A([422]), .B([424]), .Y([426]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10242 (.A([199]), .B([426]), .X([427]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10243 (.A([425]), .B([427]), .X([428]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10244 (.A([428]), .Y([429]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10245 (.A([418]), .B([429]), .Y([430]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10246 (.A([410]), .B([430]), .X([431]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10247 (.A([410]), .B([430]), .Y([432]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10248 (.A([433]), .B([417]), .Y([434]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10249 (.A([431]), .B([432]), .Y([435]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10250 (.A([39]), .B([435]), .Y([436]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10251 (.A([434]), .B([436]), .Y([437]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10252 (.A([433]), .B([438]), .Y([439]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10253 (.A([39]), .B([440]), .Y([441]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10254 (.A([439]), .B([441]), .Y([442]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10255 (.A([433]), .B([443]), .Y([444]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10256 (.A([39]), .B([445]), .Y([446]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10257 (.A([444]), .B([446]), .Y([447]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10258 (.A([433]), .B([448]), .Y([449]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10259 (.A([39]), .B([450]), .Y([451]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10260 (.A([449]), .B([451]), .Y([452]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10261 (.A([453]), .B([454]), .X([455]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10262 (.A([453]), .B([456]), .Y([457]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10263 (.A([60]), .B([454]), .Y([458]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10264 (.A([459]), .B([458]), .Y([460]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10265 (.A([457]), .B([460]), .Y([461]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10266 (.A([462]), .B([461]), .X([463]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10267 (.A([462]), .B([145]), .Y([464]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10268 (.A([463]), .B([464]), .Y([465]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10269 (.A([466]), .B([465]), .Y([467]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10270 (.A([468]), .B([469]), .X([470]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10271 (.A([470]), .Y([471]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10272 (.A([472]), .B([455]), .Y([473]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10273 (.A([474]), .B([469]), .Y([475]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10274 (.A([476]), .B([473]), .Y([477]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10275 (.A([475]), .B([477]), .X([478]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10276 (.A([467]), .B([478]), .Y([479]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10277 (.A([471]), .B([479]), .X([480]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10278 (.A([481]), .B([482]), .Y([483]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10279 (.A([484]), .B([483]), .Y([485]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10280 (.A([472]), .B([485]), .Y([486]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10281 (.A([476]), .B([486]), .Y([487]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10282 (.A([488]), .B([489]), .X([490]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10283 (.A([490]), .Y([491]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10284 (.A([469]), .B([490]), .Y([492]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10285 (.A([492]), .Y([493]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10286 (.A([494]), .B([493]), .Y([495]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10287 (.A([496]), .B([495]), .X([497]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10288 (.A([487]), .B([497]), .X([498]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10289 (.A([236]), .B([490]), .X([499]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10290 (.A([419]), .B([490]), .Y([500]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10291 (.A([501]), .B([500]), .X([502]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10292 (.A([499]), .B([502]), .Y([503]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10293 (.A([234]), .B([487]), .Y([504]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10294 (.A([492]), .B([504]), .X([505]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10295 (.A([498]), .B([505]), .Y([506]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10296 (.A([503]), .B([506]), .X([507]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10297 (.A([508]), .B([469]), .X([509]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10298 (.A([462]), .B([286]), .Y([510]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10299 (.A([511]), .B([485]), .X([512]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10300 (.A([145]), .B([169]), .X([513]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10301 (.A([191]), .B([213]), .X([514]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10302 (.A([513]), .B([514]), .X([515]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10303 (.A([234]), .B([516]), .X([517]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10304 (.A([286]), .B([518]), .X([519]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10305 (.A([517]), .B([519]), .X([520]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10306 (.A([515]), .B([520]), .X([521]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10307 (.A([462]), .B([521]), .X([522]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10308 (.A([522]), .Y([523]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10309 (.A([512]), .B([523]), .Y([524]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10310 (.A([510]), .B([524]), .Y([525]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10311 (.A([466]), .B([525]), .Y([526]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10312 (.A([509]), .B([526]), .Y([527]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10313 (.A([490]), .B([527]), .Y([528]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10314 (.A([490]), .B([521]), .X([529]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10315 (.A([472]), .B([512]), .Y([530]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10316 (.A([531]), .B([476]), .Y([532]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10317 (.A([492]), .B([532]), .X([533]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10318 (.A([533]), .Y([534]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10319 (.A([530]), .B([534]), .Y([535]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10320 (.A([529]), .B([535]), .Y([536]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10321 (.A([536]), .Y([537]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10322 (.A([528]), .B([537]), .Y([538]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10323 (.A([539]), .B([491]), .Y([540]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10324 (.A([540]), .Y([541]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10325 (.A([542]), .B([540]), .Y([543]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10326 (.A([544]), .B([539]), .X([545]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10327 (.A([546]), .B([545]), .X([547]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10328 (.A([547]), .Y([548]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10329 (.A([543]), .B([547]), .Y([549]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10330 (.A([550]), .B([549]), .X([551]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10331 (.A([60]), .B([552]), .Y([553]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10332 (.A([554]), .B([44]), .Y([555]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10333 (.A([554]), .B([553]), .X([556]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10334 (.A([555]), .B([556]), .Y([557]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10335 (.A([462]), .B([557]), .X([558]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10336 (.A([462]), .B([263]), .Y([559]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10337 (.A([558]), .B([559]), .Y([560]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10338 (.A([548]), .B([560]), .Y([561]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10339 (.A([562]), .B([472]), .Y([563]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10340 (.A([563]), .Y([564]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10341 (.A([561]), .B([564]), .Y([565]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10342 (.A([542]), .B([565]), .X([566]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10343 (.A([567]), .B([469]), .X([568]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10344 (.A([540]), .B([568]), .Y([569]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10345 (.A([569]), .Y([570]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10346 (.A([566]), .B([570]), .Y([571]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10347 (.A([551]), .B([571]), .Y([572]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10348 (.A([462]), .B([554]), .X([573]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10349 (.A([552]), .B([573]), .X([574]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10350 (.A([547]), .B([574]), .X([575]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10351 (.A([564]), .B([575]), .Y([576]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10352 (.A([577]), .B([469]), .Y([578]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10353 (.A([578]), .Y([579]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10354 (.A([576]), .B([579]), .Y([580]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10355 (.A([541]), .B([580]), .X([581]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10356 (.A([572]), .B([581]), .Y([582]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10357 (.A([433]), .B([583]), .Y([584]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10358 (.A([585]), .B([584]), .Y([586]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10359 (.A([587]), .B([588]), .X([589]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10360 (.A([590]), .B([588]), .Y([591]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10361 (.A([589]), .B([591]), .Y([592]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10362 (.A([593]), .B([592]), .Y([594]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10363 (.A([595]), .B([588]), .X([596]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10364 (.A([597]), .B([588]), .Y([598]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10365 (.A([596]), .B([598]), .Y([599]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10366 (.A([600]), .B([599]), .Y([601]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10367 (.A([594]), .B([601]), .Y([602]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10368 (.A([603]), .B([602]), .Y([604]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10369 (.A([605]), .B([606]), .X([607]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10370 (.A([608]), .B([609]), .X([610]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10371 (.A([611]), .B([610]), .X([612]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10372 (.A([607]), .B([612]), .Y([613]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10373 (.A([614]), .B([615]), .X([616]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10374 (.A([617]), .B([616]), .Y([618]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10375 (.A([613]), .B([618]), .X([619]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10376 (.A([469]), .B([150]), .Y([620]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10377 (.A([488]), .B([621]), .X([622]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10378 (.A([614]), .B([623]), .X([624]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10379 (.A([622]), .B([624]), .Y([625]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10380 (.A([620]), .B([625]), .X([626]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10381 (.A([488]), .B([623]), .X([627]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10382 (.A([627]), .Y([628]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10383 (.A([629]), .B([627]), .Y([630]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10384 (.A([605]), .B([631]), .X([632]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10385 (.A([632]), .Y([633]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10386 (.A([634]), .B([630]), .X([635]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10387 (.A([626]), .B([633]), .X([636]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10388 (.A([635]), .B([636]), .X([637]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10389 (.A([637]), .Y([638]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10390 (.A([605]), .B([639]), .X([640]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10391 (.A([641]), .B([642]), .X([643]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10392 (.A([614]), .B([643]), .X([644]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10393 (.A([640]), .B([644]), .Y([645]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10394 (.A([614]), .B([610]), .X([646]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10395 (.A([605]), .B([610]), .X([647]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10396 (.A([646]), .B([647]), .Y([648]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10397 (.A([645]), .B([648]), .X([649]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10398 (.A([650]), .B([649]), .X([651]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10399 (.A([619]), .B([651]), .X([652]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10400 (.A([637]), .B([652]), .X([653]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10401 (.A([614]), .B([654]), .X([655]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10402 (.A([655]), .Y([656]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10403 (.A([605]), .B([643]), .X([657]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10404 (.A([264]), .B([657]), .Y([658]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10405 (.A([656]), .B([658]), .X([659]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10406 (.A([488]), .B([643]), .X([660]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10407 (.A([660]), .Y([661]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10408 (.A([488]), .B([639]), .X([662]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10409 (.A([660]), .B([662]), .Y([663]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10410 (.A([491]), .B([663]), .X([664]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10411 (.A([659]), .B([664]), .X([665]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10412 (.A([666]), .B([614]), .X([667]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10413 (.A([488]), .B([606]), .X([668]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10414 (.A([667]), .B([668]), .Y([669]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10415 (.A([148]), .B([669]), .X([670]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10416 (.A([603]), .B([670]), .X([671]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10417 (.A([665]), .B([671]), .X([672]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10418 (.A([653]), .B([672]), .X([673]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10419 (.A([673]), .Y([674]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10420 (.A([675]), .B([674]), .Y([676]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10421 (.A([516]), .B([653]), .Y([677]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10422 (.A([678]), .B([665]), .Y([679]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10423 (.A([256]), .B([669]), .Y([680]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10424 (.A([681]), .B([680]), .Y([682]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10425 (.A([682]), .Y([683]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10426 (.A([679]), .B([683]), .Y([684]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10427 (.A([684]), .Y([685]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10428 (.A([677]), .B([685]), .Y([686]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10429 (.A([686]), .Y([687]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10430 (.A([676]), .B([687]), .Y([688]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10431 (.A([688]), .Y([689]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10432 (.A([604]), .B([689]), .Y([84]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10433 (.A([690]), .B([691]), .Y([692]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10434 (.A([488]), .B([610]), .X([693]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10435 (.A([694]), .B([693]), .Y([695]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10436 (.A([695]), .Y([696]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10437 (.A([697]), .B([695]), .X([698]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10438 (.A([39]), .B([692]), .Y([699]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10439 (.A([698]), .B([699]), .X([700]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10440 (.A([700]), .Y([701]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10441 (.A([84]), .B([701]), .Y([702]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10442 (.A([678]), .B([700]), .Y([703]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10443 (.A([702]), .B([703]), .Y([704]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10444 (.A([705]), .B([588]), .Y([706]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10445 (.A([707]), .B([588]), .X([708]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10446 (.A([706]), .B([708]), .Y([709]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10447 (.A([600]), .B([709]), .Y([710]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10448 (.A([711]), .B([482]), .X([712]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10449 (.A([712]), .Y([713]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10450 (.A([714]), .B([715]), .X([716]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10451 (.A([710]), .B([716]), .Y([717]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10452 (.A([713]), .B([717]), .X([718]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10453 (.A([719]), .B([718]), .X([720]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10454 (.A([721]), .B([674]), .Y([722]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10455 (.A([286]), .B([653]), .Y([723]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10456 (.A([724]), .B([665]), .Y([725]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10457 (.A([281]), .B([669]), .Y([726]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10458 (.A([725]), .B([726]), .Y([727]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10459 (.A([722]), .B([723]), .Y([728]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10460 (.A([729]), .B([728]), .X([730]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10461 (.A([727]), .B([730]), .X([731]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10462 (.A([731]), .Y([732]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10463 (.A([720]), .B([732]), .Y([85]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10464 (.A([701]), .B([85]), .Y([733]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10465 (.A([724]), .B([700]), .Y([734]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10466 (.A([733]), .B([734]), .Y([735]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10467 (.A([736]), .B([737]), .Y([738]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10468 (.A([739]), .B([588]), .Y([740]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10469 (.A([738]), .B([740]), .Y([741]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10470 (.A([593]), .B([741]), .X([742]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10471 (.A([743]), .B([482]), .X([744]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10472 (.A([744]), .Y([745]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10473 (.A([746]), .B([715]), .X([747]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10474 (.A([742]), .B([747]), .Y([748]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10475 (.A([745]), .B([748]), .X([749]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10476 (.A([719]), .B([749]), .X([750]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10477 (.A([138]), .B([674]), .Y([751]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10478 (.A([518]), .B([653]), .Y([752]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10479 (.A([753]), .B([665]), .Y([754]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10480 (.A([305]), .B([669]), .Y([755]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10481 (.A([754]), .B([755]), .Y([756]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10482 (.A([124]), .B([756]), .X([757]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10483 (.A([757]), .Y([758]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10484 (.A([752]), .B([758]), .Y([759]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10485 (.A([759]), .Y([760]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10486 (.A([751]), .B([760]), .Y([761]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10487 (.A([761]), .Y([762]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10488 (.A([750]), .B([762]), .Y([86]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10489 (.A([701]), .B([86]), .Y([763]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10490 (.A([753]), .B([700]), .Y([764]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10491 (.A([763]), .B([764]), .Y([765]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10492 (.A([766]), .B([737]), .Y([767]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10493 (.A([768]), .B([588]), .Y([769]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10494 (.A([767]), .B([769]), .Y([770]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10495 (.A([593]), .B([770]), .X([771]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10496 (.A([772]), .B([715]), .X([773]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10497 (.A([773]), .Y([774]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10498 (.A([775]), .B([482]), .X([776]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10499 (.A([771]), .B([776]), .Y([777]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10500 (.A([774]), .B([777]), .X([778]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10501 (.A([719]), .B([778]), .X([779]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10502 (.A([142]), .B([674]), .Y([780]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10503 (.A([145]), .B([653]), .Y([781]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10504 (.A([152]), .B([665]), .Y([782]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10505 (.A([329]), .B([669]), .Y([783]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10506 (.A([149]), .B([783]), .Y([784]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10507 (.A([784]), .Y([785]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10508 (.A([782]), .B([785]), .Y([786]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10509 (.A([786]), .Y([787]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10510 (.A([781]), .B([787]), .Y([788]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10511 (.A([788]), .Y([789]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10512 (.A([780]), .B([789]), .Y([790]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10513 (.A([790]), .Y([791]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10514 (.A([779]), .B([791]), .Y([87]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10515 (.A([152]), .B([700]), .Y([792]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10516 (.A([701]), .B([87]), .Y([793]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10517 (.A([792]), .B([793]), .Y([794]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10518 (.A([795]), .B([737]), .Y([796]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10519 (.A([797]), .B([588]), .Y([798]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10520 (.A([796]), .B([798]), .Y([799]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10521 (.A([593]), .B([799]), .X([800]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10522 (.A([801]), .B([482]), .X([802]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10523 (.A([802]), .Y([803]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10524 (.A([804]), .B([715]), .X([805]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10525 (.A([800]), .B([805]), .Y([806]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10526 (.A([803]), .B([806]), .X([807]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10527 (.A([719]), .B([807]), .X([808]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10528 (.A([167]), .B([674]), .Y([809]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10529 (.A([169]), .B([653]), .Y([810]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10530 (.A([175]), .B([665]), .Y([811]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10531 (.A([352]), .B([669]), .Y([812]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10532 (.A([173]), .B([812]), .Y([813]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10533 (.A([813]), .Y([814]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10534 (.A([811]), .B([814]), .Y([815]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10535 (.A([815]), .Y([816]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10536 (.A([810]), .B([816]), .Y([817]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10537 (.A([817]), .Y([818]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10538 (.A([809]), .B([818]), .Y([819]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10539 (.A([819]), .Y([820]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10540 (.A([808]), .B([820]), .Y([88]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10541 (.A([701]), .B([88]), .Y([821]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10542 (.A([175]), .B([700]), .Y([822]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10543 (.A([821]), .B([822]), .Y([823]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10544 (.A([824]), .B([737]), .Y([825]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10545 (.A([826]), .B([588]), .Y([827]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10546 (.A([825]), .B([827]), .Y([828]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10547 (.A([593]), .B([828]), .X([829]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10548 (.A([830]), .B([482]), .X([831]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10549 (.A([831]), .Y([832]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10550 (.A([833]), .B([715]), .X([834]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10551 (.A([829]), .B([834]), .Y([835]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10552 (.A([832]), .B([835]), .X([836]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10553 (.A([719]), .B([836]), .X([837]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10554 (.A([189]), .B([674]), .Y([838]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10555 (.A([191]), .B([653]), .Y([839]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10556 (.A([194]), .B([665]), .Y([840]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10557 (.A([375]), .B([669]), .Y([841]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10558 (.A([193]), .B([841]), .Y([842]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10559 (.A([842]), .Y([843]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10560 (.A([840]), .B([843]), .Y([844]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10561 (.A([844]), .Y([845]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10562 (.A([839]), .B([845]), .Y([846]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10563 (.A([846]), .Y([847]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10564 (.A([838]), .B([847]), .Y([848]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10565 (.A([848]), .Y([849]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10566 (.A([837]), .B([849]), .Y([89]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10567 (.A([701]), .B([89]), .Y([850]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10568 (.A([194]), .B([700]), .Y([851]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10569 (.A([850]), .B([851]), .Y([852]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10570 (.A([853]), .B([737]), .Y([854]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10571 (.A([855]), .B([588]), .Y([856]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10572 (.A([854]), .B([856]), .Y([857]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10573 (.A([593]), .B([857]), .X([858]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10574 (.A([859]), .B([482]), .X([860]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10575 (.A([860]), .Y([861]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10576 (.A([862]), .B([715]), .X([863]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10577 (.A([858]), .B([863]), .Y([864]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10578 (.A([861]), .B([864]), .X([865]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10579 (.A([719]), .B([865]), .X([866]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10580 (.A([211]), .B([674]), .Y([867]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10581 (.A([213]), .B([653]), .Y([868]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10582 (.A([218]), .B([665]), .Y([869]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10583 (.A([398]), .B([669]), .Y([870]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10584 (.A([216]), .B([870]), .Y([871]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10585 (.A([871]), .Y([872]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10586 (.A([869]), .B([872]), .Y([873]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10587 (.A([873]), .Y([874]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10588 (.A([868]), .B([874]), .Y([875]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10589 (.A([875]), .Y([876]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10590 (.A([867]), .B([876]), .Y([877]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10591 (.A([877]), .Y([878]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10592 (.A([866]), .B([878]), .Y([90]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10593 (.A([218]), .B([700]), .Y([879]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10594 (.A([701]), .B([90]), .Y([880]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10595 (.A([879]), .B([880]), .Y([881]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10596 (.A([882]), .B([737]), .Y([883]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10597 (.A([884]), .B([588]), .Y([885]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10598 (.A([883]), .B([885]), .Y([886]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10599 (.A([593]), .B([886]), .X([887]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10600 (.A([888]), .B([715]), .X([889]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10601 (.A([889]), .Y([890]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10602 (.A([891]), .B([482]), .X([892]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10603 (.A([887]), .B([892]), .Y([893]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10604 (.A([890]), .B([893]), .X([894]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10605 (.A([719]), .B([894]), .X([895]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10606 (.A([232]), .B([674]), .Y([896]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10607 (.A([234]), .B([653]), .Y([897]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10608 (.A([239]), .B([665]), .Y([898]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10609 (.A([419]), .B([669]), .Y([899]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10610 (.A([899]), .Y([900]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10611 (.A([237]), .B([895]), .Y([901]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10612 (.A([897]), .B([898]), .Y([902]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10613 (.A([902]), .Y([903]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10614 (.A([896]), .B([903]), .Y([904]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10615 (.A([900]), .B([904]), .X([905]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10616 (.A([901]), .B([905]), .X([91]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10617 (.A([701]), .B([91]), .Y([906]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10618 (.A([239]), .B([700]), .Y([907]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10619 (.A([906]), .B([907]), .Y([908]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10620 (.A([253]), .B([674]), .Y([909]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10621 (.A([256]), .B([651]), .Y([910]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10622 (.A([638]), .B([910]), .Y([911]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10623 (.A([719]), .B([260]), .Y([912]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10624 (.A([258]), .B([664]), .Y([913]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10625 (.A([516]), .B([659]), .Y([914]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10626 (.A([913]), .B([914]), .Y([915]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10627 (.A([912]), .B([915]), .X([916]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10628 (.A([911]), .B([916]), .X([917]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10629 (.A([917]), .Y([918]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10630 (.A([909]), .B([918]), .Y([92]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10631 (.A([258]), .B([700]), .Y([919]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10632 (.A([701]), .B([92]), .Y([920]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10633 (.A([919]), .B([920]), .Y([921]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10634 (.A([279]), .B([674]), .Y([922]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10635 (.A([281]), .B([651]), .Y([923]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10636 (.A([283]), .B([664]), .Y([924]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10637 (.A([286]), .B([659]), .Y([925]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10638 (.A([285]), .B([925]), .Y([926]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10639 (.A([923]), .B([924]), .Y([927]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10640 (.A([926]), .B([927]), .X([928]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10641 (.A([928]), .Y([929]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10642 (.A([922]), .B([929]), .Y([93]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10643 (.A([283]), .B([700]), .Y([930]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10644 (.A([701]), .B([93]), .Y([931]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10645 (.A([930]), .B([931]), .Y([932]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10646 (.A([303]), .B([674]), .Y([933]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10647 (.A([305]), .B([651]), .Y([934]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10648 (.A([518]), .B([659]), .Y([935]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10649 (.A([307]), .B([664]), .Y([936]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10650 (.A([934]), .B([936]), .Y([937]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10651 (.A([311]), .B([935]), .Y([938]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10652 (.A([937]), .B([938]), .X([939]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10653 (.A([939]), .Y([940]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10654 (.A([933]), .B([940]), .Y([94]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10655 (.A([307]), .B([700]), .Y([941]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10656 (.A([701]), .B([94]), .Y([942]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10657 (.A([941]), .B([942]), .Y([943]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10658 (.A([327]), .B([674]), .Y([944]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10659 (.A([329]), .B([651]), .Y([945]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10660 (.A([145]), .B([659]), .Y([946]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10661 (.A([331]), .B([664]), .Y([947]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10662 (.A([334]), .B([947]), .Y([948]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10663 (.A([945]), .B([946]), .Y([949]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10664 (.A([948]), .B([949]), .X([950]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10665 (.A([950]), .Y([951]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10666 (.A([944]), .B([951]), .Y([95]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10667 (.A([701]), .B([95]), .Y([952]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10668 (.A([331]), .B([700]), .Y([953]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10669 (.A([952]), .B([953]), .Y([954]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10670 (.A([349]), .B([674]), .Y([955]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10671 (.A([352]), .B([651]), .Y([956]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10672 (.A([169]), .B([659]), .Y([957]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10673 (.A([355]), .B([664]), .Y([958]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10674 (.A([956]), .B([958]), .Y([959]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10675 (.A([358]), .B([957]), .Y([960]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10676 (.A([959]), .B([960]), .X([961]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10677 (.A([961]), .Y([962]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10678 (.A([955]), .B([962]), .Y([96]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10679 (.A([701]), .B([96]), .Y([963]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10680 (.A([355]), .B([700]), .Y([964]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10681 (.A([963]), .B([964]), .Y([965]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10682 (.A([373]), .B([674]), .Y([966]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10683 (.A([375]), .B([651]), .Y([967]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10684 (.A([378]), .B([664]), .Y([968]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10685 (.A([191]), .B([659]), .Y([969]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10686 (.A([380]), .B([969]), .Y([970]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10687 (.A([967]), .B([968]), .Y([971]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10688 (.A([970]), .B([971]), .X([972]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10689 (.A([972]), .Y([973]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10690 (.A([966]), .B([973]), .Y([97]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10691 (.A([701]), .B([97]), .Y([974]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10692 (.A([378]), .B([700]), .Y([975]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10693 (.A([974]), .B([975]), .Y([976]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10694 (.A([396]), .B([674]), .Y([977]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10695 (.A([398]), .B([651]), .Y([978]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10696 (.A([978]), .Y([979]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10697 (.A([213]), .B([659]), .Y([980]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10698 (.A([980]), .Y([981]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10699 (.A([400]), .B([664]), .Y([982]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10700 (.A([401]), .B([982]), .Y([983]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10701 (.A([981]), .B([983]), .X([984]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10702 (.A([979]), .B([984]), .X([985]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10703 (.A([985]), .Y([986]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10704 (.A([977]), .B([986]), .Y([98]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10705 (.A([701]), .B([98]), .Y([987]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10706 (.A([400]), .B([700]), .Y([988]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10707 (.A([987]), .B([988]), .Y([989]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10708 (.A([417]), .B([674]), .Y([990]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10709 (.A([419]), .B([651]), .Y([991]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10710 (.A([234]), .B([659]), .Y([992]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10711 (.A([421]), .B([664]), .Y([993]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10712 (.A([424]), .B([993]), .Y([994]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10713 (.A([991]), .B([992]), .Y([995]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10714 (.A([994]), .B([995]), .X([996]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10715 (.A([996]), .Y([997]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10716 (.A([990]), .B([997]), .Y([99]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10717 (.A([701]), .B([99]), .Y([998]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10718 (.A([421]), .B([700]), .Y([999]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10719 (.A([998]), .B([999]), .Y([1000]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10720 (.A([39]), .B([695]), .Y([1001]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10721 (.A([1002]), .B([1001]), .X([1003]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10722 (.A([1003]), .Y([1004]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10723 (.A([567]), .B([1003]), .X([1005]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10724 (.A([1006]), .B([1003]), .Y([1007]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10725 (.A([1005]), .B([1007]), .Y([1008]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10726 (.A([508]), .B([1003]), .X([1009]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10727 (.A([1010]), .B([1003]), .Y([1011]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10728 (.A([1009]), .B([1011]), .Y([1012]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10729 (.A([1013]), .B([1003]), .Y([1014]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10730 (.A([1015]), .B([1003]), .X([1016]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10731 (.A([1014]), .B([1016]), .Y([1017]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10732 (.A([468]), .B([1003]), .X([1018]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10733 (.A([1019]), .B([1003]), .Y([1020]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10734 (.A([1018]), .B([1020]), .Y([1021]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10735 (.A([352]), .B([1004]), .Y([1022]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10736 (.A([1023]), .B([1003]), .Y([1024]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10737 (.A([1022]), .B([1024]), .Y([1025]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10738 (.A([1026]), .B([1003]), .Y([1027]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10739 (.A([1028]), .B([1003]), .X([1029]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10740 (.A([1027]), .B([1029]), .Y([1030]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10741 (.A([1031]), .B([1003]), .Y([1032]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10742 (.A([1033]), .B([1003]), .X([1034]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10743 (.A([1032]), .B([1034]), .Y([1035]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10744 (.A([1036]), .B([1003]), .Y([1037]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10745 (.A([419]), .B([1004]), .Y([1038]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10746 (.A([1037]), .B([1038]), .Y([1039]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10747 (.A([1040]), .B([1041]), .Y([1042]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10748 (.A([1043]), .B([1042]), .Y([1044]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10749 (.A([1044]), .Y([1045]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10750 (.A([1046]), .B([1047]), .X([1048]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10751 (.A([1049]), .B([1050]), .X([1051]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10752 (.A([1052]), .B([1051]), .X([1053]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10753 (.A([1048]), .B([1053]), .Y([1054]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10754 (.A([1055]), .B([1056]), .X([1057]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10755 (.A([1058]), .B([1057]), .X([1059]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10756 (.A([1059]), .Y([1060]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10757 (.A([1061]), .B([1062]), .X([1063]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10758 (.A([1064]), .B([1063]), .Y([1065]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10759 (.A([1066]), .B([1065]), .X([1067]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10760 (.A([1060]), .B([1067]), .X([1068]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10761 (.A([1069]), .B([1062]), .Y([1070]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10762 (.A([1070]), .Y([1071]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10763 (.A([1072]), .B([1073]), .Y([1074]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10764 (.A([1071]), .B([1074]), .Y([1075]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10765 (.A([1047]), .B([1076]), .X([1077]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10766 (.A([1077]), .Y([1078]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10767 (.A([1075]), .B([1077]), .Y([1079]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10768 (.A([1068]), .B([1079]), .X([1080]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10769 (.A([1054]), .B([1080]), .X([1081]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10770 (.A([1045]), .B([1081]), .X([1082]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10771 (.A([1083]), .B([1047]), .X([1084]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10772 (.A([1085]), .B([1084]), .Y([1086]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10773 (.A([1087]), .B([1088]), .X([1089]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10774 (.A([1057]), .B([1089]), .X([1090]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10775 (.A([1052]), .B([1089]), .X([1091]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10776 (.A([1090]), .B([1091]), .Y([1092]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10777 (.A([1086]), .B([1092]), .X([1093]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10778 (.A([1094]), .B([1095]), .X([1096]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10779 (.A([1097]), .B([1041]), .X([1098]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10780 (.A([1056]), .B([1098]), .X([1099]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10781 (.A([1096]), .B([1099]), .Y([1100]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10782 (.A([1101]), .B([1057]), .X([1102]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10783 (.A([1095]), .B([1070]), .Y([1103]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10784 (.A([1094]), .B([1103]), .Y([1104]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10785 (.A([1046]), .B([1057]), .X([1105]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10786 (.A([1104]), .B([1105]), .Y([1106]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10787 (.A([1106]), .Y([1107]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10788 (.A([1102]), .B([1107]), .Y([1108]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10789 (.A([1100]), .B([1108]), .X([1109]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10790 (.A([1093]), .B([1109]), .X([1110]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10791 (.A([1082]), .B([1110]), .X([1111]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10792 (.A([264]), .B([692]), .Y([1112]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10793 (.A([1113]), .B([660]), .Y([1114]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10794 (.A([1115]), .B([1114]), .X([1116]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10795 (.A([1112]), .B([1116]), .X([1117]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10796 (.A([646]), .B([655]), .Y([1118]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10797 (.A([1119]), .B([1118]), .X([1120]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10798 (.A([491]), .B([1120]), .X([1121]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10799 (.A([1121]), .Y([1122]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10800 (.A([1123]), .B([691]), .Y([1124]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10801 (.A([1125]), .B([1126]), .Y([1127]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10802 (.A([1127]), .Y([1128]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10803 (.A([1124]), .B([1128]), .Y([1129]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10804 (.A([617]), .B([1130]), .Y([1131]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10805 (.A([1132]), .B([1133]), .Y([1134]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10806 (.A([1131]), .B([1134]), .X([1135]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10807 (.A([1129]), .B([1135]), .X([1136]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10808 (.A([1121]), .B([1136]), .X([1137]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10809 (.A([1117]), .B([1137]), .X([1138]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10810 (.A([469]), .B([622]), .Y([1139]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10811 (.A([630]), .B([1139]), .X([1140]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10812 (.A([1141]), .B([1140]), .X([1142]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10813 (.A([1143]), .B([1144]), .X([1145]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10814 (.A([1142]), .B([1145]), .X([1146]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10815 (.A([645]), .B([695]), .X([1147]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10816 (.A([647]), .B([657]), .Y([1148]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10817 (.A([624]), .B([632]), .Y([1149]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10818 (.A([1148]), .B([1149]), .X([1150]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10819 (.A([1147]), .B([1150]), .X([1151]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10820 (.A([662]), .B([668]), .Y([1152]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10821 (.A([614]), .B([1153]), .X([1154]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10822 (.A([1154]), .Y([1155]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10823 (.A([614]), .B([621]), .X([1156]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10824 (.A([1156]), .Y([1157]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10825 (.A([1154]), .B([1156]), .Y([1158]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10826 (.A([1152]), .B([1158]), .X([1159]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10827 (.A([1160]), .B([1161]), .Y([1162]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10828 (.A([613]), .B([1162]), .X([1163]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10829 (.A([1159]), .B([1163]), .X([1164]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10830 (.A([1151]), .B([1164]), .X([1165]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10831 (.A([1146]), .B([1165]), .X([1166]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10832 (.A([1138]), .B([1166]), .X([1167]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10833 (.A([39]), .B([1167]), .Y([1168]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10834 (.A([1168]), .Y([1169]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10835 (.A([1051]), .B([1057]), .X([1170]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10836 (.A([1040]), .B([1057]), .X([1171]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10837 (.A([1111]), .B([1169]), .Y([1172]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10838 (.A([1172]), .Y([1173]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10839 (.A([1174]), .B([1063]), .X([1175]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10840 (.A([1175]), .Y([1176]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10841 (.A([1100]), .B([1176]), .X([1177]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10842 (.A([1060]), .B([1177]), .X([1178]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10843 (.A([1077]), .B([1090]), .Y([1179]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10844 (.A([1178]), .B([1179]), .X([1180]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10845 (.A([472]), .B([1180]), .Y([1181]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10846 (.A([612]), .B([668]), .Y([1182]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10847 (.A([1148]), .B([1182]), .X([1183]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10848 (.A([172]), .B([1184]), .X([1185]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10849 (.A([1156]), .B([1185]), .Y([1186]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10850 (.A([1160]), .B([150]), .Y([1187]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10851 (.A([1161]), .B([1188]), .Y([1189]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10852 (.A([1187]), .B([1189]), .X([1190]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10853 (.A([1186]), .B([1190]), .X([1191]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10854 (.A([1183]), .B([1191]), .X([1192]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10855 (.A([1193]), .B([550]), .X([1194]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10856 (.A([1194]), .Y([1195]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10857 (.A([1196]), .B([1194]), .X([1197]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10858 (.A([640]), .B([1197]), .X([1198]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10859 (.A([1124]), .B([1198]), .Y([1199]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10860 (.A([1200]), .B([1201]), .Y([1202]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10861 (.A([1199]), .B([1202]), .X([1203]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10862 (.A([1130]), .B([622]), .Y([1204]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10863 (.A([1155]), .B([1204]), .X([1205]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10864 (.A([629]), .B([694]), .Y([1206]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10865 (.A([1133]), .B([644]), .Y([1207]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10866 (.A([1206]), .B([1207]), .X([1208]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10867 (.A([1205]), .B([1208]), .X([1209]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10868 (.A([1203]), .B([1209]), .X([1210]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10869 (.A([1121]), .B([1210]), .X([1211]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10870 (.A([1192]), .B([1211]), .X([1212]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10871 (.A([1212]), .Y([1213]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10872 (.A([1181]), .B([1213]), .Y([1214]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10873 (.A([1173]), .B([1214]), .Y([1215]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10874 (.A([1216]), .B([1172]), .Y([1217]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10875 (.A([1215]), .B([1217]), .Y([1218]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10876 (.A([1219]), .B([1091]), .Y([1220]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10877 (.A([1094]), .B([1064]), .X([1221]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10878 (.A([1048]), .B([1221]), .Y([1222]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10879 (.A([1222]), .Y([1223]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10880 (.A([1106]), .B([1176]), .X([1224]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10881 (.A([1222]), .B([1224]), .X([1225]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10882 (.A([1220]), .B([1225]), .X([1226]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10883 (.A([472]), .B([1226]), .Y([1227]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10884 (.A([438]), .B([443]), .X([1228]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10885 (.A([1228]), .Y([1229]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10886 (.A([1230]), .B([1229]), .Y([1231]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10887 (.A([438]), .B([1232]), .X([1233]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10888 (.A([1233]), .Y([1234]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10889 (.A([1235]), .B([1234]), .Y([1236]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10890 (.A([1231]), .B([1236]), .Y([1237]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10891 (.A([1238]), .B([1232]), .X([1239]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10892 (.A([1240]), .B([1239]), .X([1241]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10893 (.A([443]), .B([1238]), .X([1242]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10894 (.A([1243]), .B([1242]), .X([1244]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10895 (.A([1241]), .B([1244]), .Y([1245]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10896 (.A([1237]), .B([1245]), .X([1246]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10897 (.A([1247]), .B([1246]), .Y([1248]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10898 (.A([1249]), .B([1229]), .Y([1250]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10899 (.A([1251]), .B([1234]), .Y([1252]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10900 (.A([1250]), .B([1252]), .Y([1253]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10901 (.A([1254]), .B([1239]), .X([1255]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10902 (.A([496]), .B([1242]), .X([1256]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10903 (.A([1255]), .B([1256]), .Y([1257]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10904 (.A([1253]), .B([1257]), .X([1258]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10905 (.A([1259]), .B([1258]), .Y([1260]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10906 (.A([1248]), .B([1260]), .Y([1261]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10907 (.A([1262]), .B([1261]), .Y([1263]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10908 (.A([1264]), .B([1265]), .X([1266]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10909 (.A([1266]), .Y([1267]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10910 (.A([622]), .B([667]), .Y([1268]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10911 (.A([633]), .B([1268]), .X([1269]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10912 (.A([1186]), .B([1269]), .X([1270]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10913 (.A([1266]), .B([1270]), .X([1271]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10914 (.A([1196]), .B([1183]), .Y([1272]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10915 (.A([1272]), .Y([1273]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10916 (.A([1274]), .B([150]), .Y([1275]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10917 (.A([1276]), .B([1275]), .X([1277]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10918 (.A([662]), .B([693]), .Y([1278]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10919 (.A([1127]), .B([1278]), .X([1279]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10920 (.A([1277]), .B([1279]), .X([1280]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10921 (.A([1280]), .Y([1281]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10922 (.A([1263]), .B([1281]), .Y([1282]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10923 (.A([1271]), .B([1282]), .X([1283]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10924 (.A([1273]), .B([1283]), .X([1284]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10925 (.A([1284]), .Y([1285]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10926 (.A([1227]), .B([1285]), .Y([1286]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10927 (.A([1172]), .B([1286]), .X([1287]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10928 (.A([1288]), .B([1173]), .X([1289]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10929 (.A([1287]), .B([1289]), .Y([1290]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10930 (.A([1290]), .Y([1291]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10931 (.A([1178]), .B([1222]), .X([1292]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10932 (.A([1093]), .B([1292]), .X([1293]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10933 (.A([472]), .B([1293]), .Y([1294]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10934 (.A([172]), .B([1295]), .Y([1296]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10935 (.A([625]), .B([1296]), .X([1297]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10936 (.A([645]), .B([1157]), .X([1298]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10937 (.A([630]), .B([1127]), .X([1299]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10938 (.A([1298]), .B([1299]), .X([1300]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10939 (.A([1297]), .B([1300]), .X([1301]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10940 (.A([1132]), .B([1302]), .Y([1303]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10941 (.A([694]), .B([662]), .Y([1304]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10942 (.A([1304]), .Y([1305]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10943 (.A([1131]), .B([1304]), .X([1306]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10944 (.A([1303]), .B([1306]), .X([1307]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10945 (.A([1117]), .B([1307]), .X([1308]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10946 (.A([1301]), .B([1308]), .X([1309]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10947 (.A([562]), .B([1183]), .Y([1310]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10948 (.A([1122]), .B([1310]), .Y([1311]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10949 (.A([1311]), .Y([1312]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10950 (.A([1294]), .B([1312]), .Y([1313]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10951 (.A([1309]), .B([1313]), .X([1314]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10952 (.A([1173]), .B([1314]), .Y([1315]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10953 (.A([1316]), .B([1172]), .Y([1317]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10954 (.A([1315]), .B([1317]), .Y([1318]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10955 (.A([1053]), .B([1105]), .Y([1319]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10956 (.A([1102]), .B([1223]), .Y([1320]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10957 (.A([1319]), .B([1320]), .X([1321]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10958 (.A([1177]), .B([1321]), .X([1322]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10959 (.A([472]), .B([1322]), .Y([1323]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10960 (.A([644]), .B([1194]), .X([1324]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10961 (.A([1324]), .Y([1325]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10962 (.A([1198]), .B([1305]), .Y([1326]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10963 (.A([1325]), .B([1326]), .X([1327]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10964 (.A([1117]), .B([1327]), .X([1328]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10965 (.A([1130]), .B([469]), .Y([1329]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10966 (.A([1329]), .Y([1330]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10967 (.A([1331]), .B([1330]), .Y([1332]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10968 (.A([630]), .B([1149]), .X([1333]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10969 (.A([1332]), .B([1333]), .X([1334]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10970 (.A([1335]), .B([1155]), .X([1336]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10971 (.A([1190]), .B([1336]), .X([1337]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10972 (.A([1334]), .B([1337]), .X([1338]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10973 (.A([1328]), .B([1338]), .X([1339]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10974 (.A([1295]), .B([1261]), .X([1340]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10975 (.A([1312]), .B([1340]), .Y([1341]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10976 (.A([1339]), .B([1341]), .X([1342]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10977 (.A([1342]), .Y([1343]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10978 (.A([1323]), .B([1343]), .Y([1344]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10979 (.A([1173]), .B([1344]), .Y([1345]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10980 (.A([1346]), .B([1172]), .Y([1347]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10981 (.A([1345]), .B([1347]), .Y([1348]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10982 (.A([1349]), .B([1063]), .X([1350]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10983 (.A([1171]), .B([1350]), .Y([1351]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10984 (.A([1054]), .B([1351]), .X([1352]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10985 (.A([1220]), .B([1352]), .X([1353]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10986 (.A([472]), .B([1353]), .Y([1354]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10987 (.A([644]), .B([1195]), .X([1355]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10988 (.A([694]), .B([607]), .Y([1356]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10989 (.A([624]), .B([1156]), .Y([1357]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10990 (.A([1356]), .B([1357]), .X([1358]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10991 (.A([1359]), .B([1127]), .X([1360]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10992 (.A([1358]), .B([1360]), .X([1361]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10993 (.A([1336]), .B([1361]), .X([1362]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10994 (.A([1124]), .B([1355]), .Y([1363]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10995 (.A([1363]), .Y([1364]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10996 (.A([1354]), .B([1364]), .Y([1365]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10997 (.A([1362]), .B([1365]), .X([1366]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10998 (.A([1173]), .B([1366]), .Y([1367]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10999 (.A([1368]), .B([1172]), .Y([1369]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11000 (.A([1367]), .B([1369]), .Y([1370]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11001 (.A([1063]), .B([1170]), .Y([1371]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11002 (.A([1086]), .B([1179]), .X([1372]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11003 (.A([1371]), .B([1372]), .X([1373]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11004 (.A([472]), .B([1373]), .Y([1374]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11005 (.A([1134]), .B([1189]), .X([1375]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11006 (.A([697]), .B([1278]), .X([1376]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11007 (.A([1273]), .B([1376]), .X([1377]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11008 (.A([1375]), .B([1377]), .X([1378]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11009 (.A([1378]), .Y([1379]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11010 (.A([1374]), .B([1379]), .Y([1380]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11011 (.A([1140]), .B([1380]), .X([1381]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11012 (.A([1173]), .B([1381]), .Y([1382]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11013 (.A([1383]), .B([1172]), .Y([1384]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11014 (.A([1382]), .B([1384]), .Y([1385]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11015 (.A([1386]), .B([1387]), .X([1388]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11016 (.A([1047]), .B([1389]), .X([1390]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11017 (.A([1349]), .B([1069]), .X([1391]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11018 (.A([1391]), .Y([1392]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11019 (.A([1049]), .B([1393]), .X([1394]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11020 (.A([1395]), .B([1394]), .X([1396]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11021 (.A([1072]), .B([1397]), .X([1398]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11022 (.A([1055]), .B([1397]), .X([1399]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11023 (.A([1392]), .B([1399]), .X([1400]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11024 (.A([1390]), .B([1400]), .Y([1401]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11025 (.A([1396]), .B([1398]), .Y([1402]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11026 (.A([1401]), .B([1402]), .X([1403]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11027 (.A([1404]), .B([1403]), .X([1405]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11028 (.A([1406]), .B([1405]), .X([1407]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11029 (.A([1388]), .B([1407]), .Y([1408]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11030 (.A([1408]), .Y([1409]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11031 (.A([1410]), .B([1387]), .X([1411]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11032 (.A([1412]), .B([1413]), .X([1414]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11033 (.A([1085]), .B([1414]), .X([1415]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11034 (.A([1415]), .Y([1416]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11035 (.A([1078]), .B([1401]), .X([1417]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11036 (.A([1416]), .B([1417]), .X([1418]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11037 (.A([1404]), .B([1418]), .X([1419]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11038 (.A([1411]), .B([1419]), .Y([1420]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11039 (.A([1420]), .Y([1421]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11040 (.A([1422]), .B([1404]), .Y([1423]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11041 (.A([1395]), .B([1414]), .X([1424]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11042 (.A([1061]), .B([440]), .X([1425]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11043 (.A([1413]), .B([1425]), .X([1426]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11044 (.A([1426]), .Y([1427]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11045 (.A([1428]), .B([1424]), .Y([1429]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11046 (.A([1427]), .B([1429]), .X([1430]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11047 (.A([1431]), .B([1430]), .Y([1432]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11048 (.A([1387]), .B([1390]), .Y([1433]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11049 (.A([1433]), .Y([1434]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11050 (.A([1432]), .B([1434]), .Y([1435]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11051 (.A([1436]), .B([1425]), .Y([1437]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11052 (.A([1438]), .B([1437]), .Y([1439]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11053 (.A([1394]), .B([1439]), .Y([1440]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11054 (.A([1406]), .B([1440]), .X([1441]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11055 (.A([1435]), .B([1441]), .X([1442]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11056 (.A([1423]), .B([1442]), .Y([1443]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11057 (.A([1443]), .Y([1444]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11058 (.A([1085]), .B([1445]), .X([1446]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11059 (.A([1446]), .Y([1447]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11060 (.A([1435]), .B([1447]), .X([1448]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11061 (.A([1449]), .B([1387]), .X([1450]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11062 (.A([1448]), .B([1450]), .Y([1451]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11063 (.A([1451]), .Y([1452]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11064 (.A([1453]), .B([1387]), .X([1454]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11065 (.A([1455]), .B([1456]), .Y([1457]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11066 (.A([1073]), .B([1457]), .X([1458]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11067 (.A([1458]), .Y([1459]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11068 (.A([1460]), .B([1072]), .X([1461]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11069 (.A([1461]), .Y([1462]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11070 (.A([1463]), .B([1464]), .Y([1465]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11071 (.A([1462]), .B([1465]), .X([1466]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11072 (.A([1404]), .B([1466]), .X([1467]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11073 (.A([1459]), .B([1465]), .X([1468]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11074 (.A([1468]), .Y([1469]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11075 (.A([1459]), .B([1467]), .X([1470]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11076 (.A([1454]), .B([1470]), .Y([1471]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11077 (.A([1471]), .Y([1472]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11078 (.A([440]), .B([1473]), .X([1474]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11079 (.A([1474]), .Y([1475]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11080 (.A([445]), .B([1390]), .X([1476]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11081 (.A([1477]), .B([1073]), .X([1478]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11082 (.A([1479]), .B([1478]), .Y([1480]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11083 (.A([1480]), .Y([1481]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11084 (.A([1476]), .B([1481]), .Y([1482]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11085 (.A([1475]), .B([1482]), .X([1483]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11086 (.A([1484]), .B([1483]), .X([1485]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11087 (.A([1468]), .B([1485]), .X([1486]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11088 (.A([1387]), .B([1486]), .Y([1487]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11089 (.A([1488]), .B([1404]), .Y([1489]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11090 (.A([1487]), .B([1489]), .Y([1490]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11091 (.A([1491]), .B([1387]), .X([1492]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11092 (.A([1462]), .B([1486]), .X([1493]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11093 (.A([1387]), .B([1493]), .Y([1494]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11094 (.A([1072]), .B([1495]), .Y([1496]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11095 (.A([1497]), .B([1496]), .Y([1498]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11096 (.A([1498]), .Y([1499]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11097 (.A([1485]), .B([1499]), .X([1500]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11098 (.A([1494]), .B([1500]), .X([1501]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11099 (.A([1492]), .B([1501]), .Y([1502]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11100 (.A([1502]), .Y([1503]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11101 (.A([1504]), .B([1387]), .X([1505]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11102 (.A([1506]), .B([1458]), .X([1507]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11103 (.A([1507]), .Y([1508]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11104 (.A([1467]), .B([1508]), .X([1509]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11105 (.A([1469]), .B([1509]), .X([1510]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11106 (.A([1505]), .B([1510]), .Y([1511]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11107 (.A([1511]), .Y([1512]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11108 (.A([433]), .B([1513]), .Y([1514]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11109 (.A([148]), .B([645]), .X([1515]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11110 (.A([1066]), .B([647]), .Y([1516]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11111 (.A([1517]), .B([663]), .X([1518]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11112 (.A([456]), .B([1518]), .X([1519]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11113 (.A([1516]), .B([1519]), .X([1520]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11114 (.A([1515]), .B([1520]), .X([1521]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11115 (.A([1521]), .Y([1522]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11116 (.A([1523]), .B([577]), .Y([1524]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11117 (.A([539]), .B([1525]), .X([1526]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11118 (.A([44]), .B([1526]), .Y([1527]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11119 (.A([1243]), .B([1526]), .X([1528]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11120 (.A([1527]), .B([1528]), .Y([1529]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11121 (.A([544]), .B([1529]), .X([1530]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11122 (.A([1531]), .B([544]), .Y([1532]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11123 (.A([1530]), .B([1532]), .Y([1533]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11124 (.A([1523]), .B([1533]), .X([1534]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11125 (.A([1524]), .B([1534]), .Y([1535]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11126 (.A([1517]), .B([1535]), .Y([1536]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11127 (.A([1536]), .Y([1537]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11128 (.A([550]), .B([1515]), .Y([1538]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11129 (.A([1538]), .Y([1539]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11130 (.A([607]), .B([667]), .Y([1540]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11131 (.A([628]), .B([1540]), .X([1541]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11132 (.A([1139]), .B([1541]), .X([1542]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11133 (.A([539]), .B([1543]), .X([1544]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11134 (.A([539]), .B([456]), .Y([1545]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11135 (.A([1544]), .B([1545]), .Y([1546]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11136 (.A([1523]), .B([1546]), .X([1547]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11137 (.A([1524]), .B([1547]), .Y([1548]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11138 (.A([663]), .B([1548]), .Y([1549]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11139 (.A([1267]), .B([1549]), .Y([1550]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11140 (.A([1542]), .B([1550]), .X([1551]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11141 (.A([1539]), .B([1551]), .X([1552]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11142 (.A([1537]), .B([1552]), .X([1553]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11143 (.A([1522]), .B([1553]), .X([1554]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11144 (.A([1555]), .B([1518]), .Y([1556]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11145 (.A([1519]), .B([1556]), .Y([1557]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11146 (.A([1557]), .Y([1558]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11147 (.A([1554]), .B([1558]), .X([1559]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11148 (.A([1274]), .B([1161]), .Y([1560]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11149 (.A([661]), .B([1560]), .X([1561]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11150 (.A([695]), .B([1561]), .X([1562]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11151 (.A([1563]), .B([1303]), .X([1564]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11152 (.A([1565]), .B([1564]), .X([1566]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11153 (.A([1562]), .B([1566]), .X([1567]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11154 (.A([1525]), .B([1113]), .X([1568]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11155 (.A([1568]), .Y([1569]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11156 (.A([1567]), .B([1569]), .X([1570]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11157 (.A([1570]), .Y([1571]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11158 (.A([894]), .B([1571]), .X([1572]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11159 (.A([607]), .B([632]), .Y([1573]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11160 (.A([628]), .B([1573]), .X([1574]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11161 (.A([626]), .B([1574]), .X([1575]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11162 (.A([1517]), .B([1516]), .X([1576]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11163 (.A([1295]), .B([662]), .Y([1577]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11164 (.A([1578]), .B([1577]), .X([1579]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11165 (.A([1576]), .B([1579]), .X([1580]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11166 (.A([1575]), .B([1580]), .X([1581]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11167 (.A([1567]), .B([1581]), .X([1582]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11168 (.A([1582]), .Y([1583]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11169 (.A([1525]), .B([44]), .Y([1584]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11170 (.A([1113]), .B([1584]), .X([1585]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11171 (.A([1582]), .B([1585]), .Y([1586]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11172 (.A([234]), .B([1575]), .Y([1587]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11173 (.A([419]), .B([1577]), .Y([1588]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11174 (.A([424]), .B([1588]), .Y([1589]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11175 (.A([1589]), .Y([1590]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11176 (.A([1587]), .B([1590]), .Y([1591]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11177 (.A([1586]), .B([1591]), .X([1592]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11178 (.A([1592]), .Y([1593]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11179 (.A([1572]), .B([1593]), .Y([1594]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11180 (.A([1504]), .B([1518]), .Y([1595]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11181 (.A([1595]), .Y([1596]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11182 (.A([1491]), .B([1518]), .Y([1597]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11183 (.A([1597]), .Y([1598]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11184 (.A([1599]), .B([1187]), .X([1600]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11185 (.A([1149]), .B([1600]), .X([1601]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11186 (.A([148]), .B([1601]), .X([1602]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11187 (.A([1531]), .B([663]), .X([1603]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11188 (.A([1576]), .B([1603]), .X([1604]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11189 (.A([1604]), .Y([1605]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11190 (.A([1602]), .B([1605]), .X([1606]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11191 (.A([1598]), .B([1606]), .X([1607]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11192 (.A([1596]), .B([1606]), .X([1608]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11193 (.A([1596]), .B([1607]), .X([1609]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11194 (.A([627]), .B([662]), .Y([1610]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11195 (.A([620]), .B([1610]), .X([1611]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11196 (.A([1516]), .B([1573]), .X([1612]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11197 (.A([1611]), .B([1612]), .X([1613]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11198 (.A([1297]), .B([1564]), .X([1614]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11199 (.A([1613]), .B([1614]), .X([1615]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11200 (.A([1562]), .B([1615]), .X([1616]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11201 (.A([1616]), .Y([1617]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11202 (.A([419]), .B([1617]), .Y([1618]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11203 (.A([232]), .B([1262]), .Y([1619]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11204 (.A([1618]), .B([1619]), .Y([1620]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11205 (.A([1620]), .Y([1621]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11206 (.A([1608]), .B([1621]), .X([1622]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11207 (.A([1607]), .B([1620]), .X([1623]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11208 (.A([1622]), .B([1623]), .Y([1624]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11209 (.A([1609]), .B([1624]), .Y([1625]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11210 (.A([1594]), .B([1622]), .X([1626]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11211 (.A([1626]), .Y([1627]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11212 (.A([1594]), .B([1625]), .Y([1628]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11213 (.A([1558]), .B([1628]), .Y([1629]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11214 (.A([1627]), .B([1629]), .X([1630]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11215 (.A([1559]), .B([1630]), .Y([1631]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11216 (.A([1520]), .B([1602]), .X([1632]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11217 (.A([1453]), .B([1518]), .Y([1633]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11218 (.A([1632]), .B([1633]), .Y([1634]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11219 (.A([583]), .B([148]), .Y([1635]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11220 (.A([1488]), .B([1518]), .Y([1636]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11221 (.A([1635]), .B([1636]), .Y([1637]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11222 (.A([1601]), .B([1637]), .X([1638]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11223 (.A([1638]), .Y([1639]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11224 (.A([1632]), .B([1639]), .Y([1640]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11225 (.A([1634]), .B([1638]), .X([1641]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11226 (.A([1620]), .B([1641]), .Y([1642]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11227 (.A([1634]), .B([1639]), .X([1643]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11228 (.A([1621]), .B([1643]), .Y([1644]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11229 (.A([1642]), .B([1644]), .Y([1645]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11230 (.A([1631]), .B([1645]), .Y([1646]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11231 (.A([1633]), .B([1640]), .X([1647]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11232 (.A([1647]), .Y([1648]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11233 (.A([1645]), .B([1647]), .Y([1649]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11234 (.A([1649]), .Y([1650]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11235 (.A([1646]), .B([1649]), .Y([1651]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11236 (.A([433]), .B([1651]), .X([1652]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11237 (.A([1514]), .B([1652]), .Y([1653]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11238 (.A([39]), .B([234]), .X([1654]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11239 (.A([1033]), .B([1616]), .X([1655]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11240 (.A([211]), .B([1262]), .Y([1656]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11241 (.A([1655]), .B([1656]), .Y([1657]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11242 (.A([1657]), .Y([1658]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11243 (.A([1643]), .B([1657]), .X([1659]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11244 (.A([1641]), .B([1658]), .X([1660]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11245 (.A([1659]), .B([1660]), .Y([1661]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11246 (.A([1648]), .B([1661]), .X([1662]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11247 (.A([865]), .B([1571]), .X([1663]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11248 (.A([213]), .B([1575]), .Y([1664]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11249 (.A([398]), .B([1577]), .Y([1665]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11250 (.A([401]), .B([1665]), .Y([1666]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11251 (.A([1585]), .B([1664]), .Y([1667]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11252 (.A([1583]), .B([1667]), .X([1668]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11253 (.A([1666]), .B([1668]), .X([1669]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11254 (.A([1669]), .Y([1670]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11255 (.A([1663]), .B([1670]), .Y([1671]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11256 (.A([1671]), .Y([1672]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11257 (.A([1608]), .B([1658]), .X([1673]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11258 (.A([1672]), .B([1673]), .Y([1674]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11259 (.A([1674]), .Y([1675]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11260 (.A([1607]), .B([1657]), .X([1676]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11261 (.A([1673]), .B([1676]), .Y([1677]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11262 (.A([1609]), .B([1677]), .Y([1678]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11263 (.A([1672]), .B([1678]), .X([1679]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11264 (.A([1557]), .B([1594]), .Y([1680]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11265 (.A([1558]), .B([1679]), .Y([1681]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11266 (.A([1675]), .B([1681]), .X([1682]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11267 (.A([1680]), .B([1682]), .Y([1683]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11268 (.A([1662]), .B([1683]), .Y([1684]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11269 (.A([1028]), .B([1616]), .X([1685]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11270 (.A([189]), .B([1262]), .Y([1686]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11271 (.A([1685]), .B([1686]), .Y([1687]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11272 (.A([1687]), .Y([1688]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11273 (.A([1641]), .B([1687]), .Y([1689]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11274 (.A([1643]), .B([1688]), .Y([1690]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11275 (.A([1689]), .B([1690]), .Y([1691]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11276 (.A([1647]), .B([1691]), .Y([1692]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11277 (.A([1692]), .Y([1693]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11278 (.A([836]), .B([1571]), .X([1694]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11279 (.A([191]), .B([1575]), .Y([1695]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11280 (.A([375]), .B([1577]), .Y([1696]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11281 (.A([380]), .B([1696]), .Y([1697]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11282 (.A([1697]), .Y([1698]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11283 (.A([1695]), .B([1698]), .Y([1699]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11284 (.A([1586]), .B([1699]), .X([1700]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11285 (.A([1700]), .Y([1701]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11286 (.A([1694]), .B([1701]), .Y([1702]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11287 (.A([1608]), .B([1688]), .X([1703]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11288 (.A([1607]), .B([1687]), .X([1704]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11289 (.A([1703]), .B([1704]), .Y([1705]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11290 (.A([1609]), .B([1705]), .Y([1706]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11291 (.A([1702]), .B([1703]), .X([1707]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11292 (.A([1702]), .B([1706]), .Y([1708]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11293 (.A([1707]), .B([1708]), .Y([1709]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11294 (.A([1557]), .B([1709]), .X([1710]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11295 (.A([1558]), .B([1671]), .X([1711]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11296 (.A([1710]), .B([1711]), .Y([1712]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11297 (.A([1693]), .B([1712]), .X([1713]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11298 (.A([352]), .B([1617]), .Y([1714]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11299 (.A([167]), .B([1262]), .Y([1715]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11300 (.A([1714]), .B([1715]), .Y([1716]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11301 (.A([1716]), .Y([1717]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11302 (.A([1643]), .B([1716]), .X([1718]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11303 (.A([1641]), .B([1717]), .X([1719]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11304 (.A([1718]), .B([1719]), .Y([1720]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11305 (.A([1648]), .B([1720]), .X([1721]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11306 (.A([807]), .B([1571]), .X([1722]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11307 (.A([169]), .B([1575]), .Y([1723]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11308 (.A([352]), .B([1577]), .Y([1724]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11309 (.A([358]), .B([1724]), .Y([1725]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11310 (.A([1725]), .Y([1726]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11311 (.A([1723]), .B([1726]), .Y([1727]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11312 (.A([1586]), .B([1727]), .X([1728]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11313 (.A([1728]), .Y([1729]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11314 (.A([1722]), .B([1729]), .Y([1730]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11315 (.A([1608]), .B([1717]), .X([1731]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11316 (.A([1731]), .Y([1732]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11317 (.A([1607]), .B([1716]), .X([1733]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11318 (.A([1731]), .B([1733]), .Y([1734]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11319 (.A([1609]), .B([1734]), .Y([1735]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11320 (.A([1735]), .Y([1736]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11321 (.A([1730]), .B([1736]), .Y([1737]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11322 (.A([1730]), .B([1732]), .X([1738]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11323 (.A([1738]), .Y([1739]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11324 (.A([1557]), .B([1702]), .Y([1740]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11325 (.A([1558]), .B([1737]), .Y([1741]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11326 (.A([1739]), .B([1741]), .X([1742]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11327 (.A([1740]), .B([1742]), .Y([1743]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11328 (.A([1721]), .B([1743]), .Y([1744]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11329 (.A([468]), .B([1616]), .X([1745]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11330 (.A([142]), .B([1262]), .Y([1746]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11331 (.A([1745]), .B([1746]), .Y([1747]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11332 (.A([1747]), .Y([1748]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11333 (.A([1641]), .B([1747]), .Y([1749]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11334 (.A([1643]), .B([1748]), .Y([1750]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11335 (.A([1749]), .B([1750]), .Y([1751]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11336 (.A([1647]), .B([1751]), .Y([1752]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11337 (.A([1752]), .Y([1753]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11338 (.A([778]), .B([1571]), .X([1754]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11339 (.A([145]), .B([1575]), .Y([1755]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11340 (.A([329]), .B([1577]), .Y([1756]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11341 (.A([334]), .B([1756]), .Y([1757]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11342 (.A([1757]), .Y([1758]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11343 (.A([1755]), .B([1758]), .Y([1759]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11344 (.A([1586]), .B([1759]), .X([1760]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11345 (.A([1760]), .Y([1761]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11346 (.A([1754]), .B([1761]), .Y([1762]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11347 (.A([1608]), .B([1748]), .X([1763]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11348 (.A([1607]), .B([1747]), .X([1764]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11349 (.A([1763]), .B([1764]), .Y([1765]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11350 (.A([1609]), .B([1765]), .Y([1766]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11351 (.A([1762]), .B([1763]), .X([1767]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11352 (.A([1762]), .B([1766]), .Y([1768]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11353 (.A([1767]), .B([1768]), .Y([1769]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11354 (.A([1557]), .B([1769]), .X([1770]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11355 (.A([1558]), .B([1730]), .X([1771]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11356 (.A([1770]), .B([1771]), .Y([1772]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11357 (.A([1753]), .B([1772]), .X([1773]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11358 (.A([1751]), .B([1772]), .Y([1774]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11359 (.A([1773]), .B([1774]), .Y([1775]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11360 (.A([1775]), .Y([1776]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11361 (.A([1015]), .B([1616]), .X([1777]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11362 (.A([138]), .B([1262]), .Y([1778]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11363 (.A([1777]), .B([1778]), .Y([1779]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11364 (.A([1779]), .Y([1780]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11365 (.A([1641]), .B([1779]), .Y([1781]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11366 (.A([1643]), .B([1780]), .Y([1782]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11367 (.A([1781]), .B([1782]), .Y([1783]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11368 (.A([1647]), .B([1783]), .Y([1784]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11369 (.A([1784]), .Y([1785]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11370 (.A([749]), .B([1571]), .X([1786]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11371 (.A([518]), .B([1575]), .Y([1787]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11372 (.A([305]), .B([1577]), .Y([1788]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11373 (.A([1585]), .B([1788]), .Y([1789]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11374 (.A([312]), .B([1789]), .X([1790]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11375 (.A([1790]), .Y([1791]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11376 (.A([1787]), .B([1791]), .Y([1792]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11377 (.A([1583]), .B([1792]), .X([1793]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11378 (.A([1793]), .Y([1794]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11379 (.A([1786]), .B([1794]), .Y([1795]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11380 (.A([1608]), .B([1780]), .X([1796]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11381 (.A([1607]), .B([1779]), .X([1797]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11382 (.A([1796]), .B([1797]), .Y([1798]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11383 (.A([1609]), .B([1798]), .Y([1799]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11384 (.A([1795]), .B([1796]), .X([1800]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11385 (.A([1795]), .B([1799]), .Y([1801]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11386 (.A([1800]), .B([1801]), .Y([1802]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11387 (.A([1557]), .B([1802]), .X([1803]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11388 (.A([1558]), .B([1762]), .X([1804]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11389 (.A([1803]), .B([1804]), .Y([1805]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11390 (.A([1785]), .B([1805]), .X([1806]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11391 (.A([508]), .B([1616]), .X([1807]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11392 (.A([721]), .B([1262]), .Y([1808]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11393 (.A([1807]), .B([1808]), .Y([1809]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11394 (.A([1809]), .Y([1810]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11395 (.A([1643]), .B([1809]), .X([1811]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11396 (.A([1641]), .B([1810]), .X([1812]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11397 (.A([1811]), .B([1812]), .Y([1813]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11398 (.A([1648]), .B([1813]), .X([1814]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11399 (.A([718]), .B([1571]), .X([1815]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11400 (.A([286]), .B([1575]), .Y([1816]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11401 (.A([281]), .B([1577]), .Y([1817]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11402 (.A([285]), .B([1582]), .Y([1818]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11403 (.A([1585]), .B([1817]), .Y([1819]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11404 (.A([1819]), .Y([1820]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11405 (.A([1816]), .B([1820]), .Y([1821]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11406 (.A([1818]), .B([1821]), .X([1822]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11407 (.A([1822]), .Y([1823]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11408 (.A([1815]), .B([1823]), .Y([1824]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11409 (.A([1608]), .B([1810]), .X([1825]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11410 (.A([1607]), .B([1809]), .X([1826]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11411 (.A([1825]), .B([1826]), .Y([1827]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11412 (.A([1609]), .B([1827]), .Y([1828]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11413 (.A([1824]), .B([1828]), .Y([1829]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11414 (.A([1824]), .B([1825]), .X([1830]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11415 (.A([1829]), .B([1830]), .Y([1831]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11416 (.A([1558]), .B([1831]), .Y([1832]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11417 (.A([1557]), .B([1795]), .Y([1833]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11418 (.A([1832]), .B([1833]), .Y([1834]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11419 (.A([1814]), .B([1834]), .Y([1835]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11420 (.A([567]), .B([1616]), .X([1836]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11421 (.A([675]), .B([1262]), .Y([1837]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11422 (.A([1836]), .B([1837]), .Y([1838]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11423 (.A([1838]), .Y([1839]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11424 (.A([1643]), .B([1838]), .X([1840]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11425 (.A([1641]), .B([1839]), .X([1841]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11426 (.A([1840]), .B([1841]), .Y([1842]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11427 (.A([1648]), .B([1842]), .X([1843]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11428 (.A([1557]), .B([1824]), .Y([1844]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11429 (.A([602]), .B([1570]), .Y([1845]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11430 (.A([516]), .B([1575]), .Y([1846]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11431 (.A([256]), .B([1577]), .Y([1847]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11432 (.A([260]), .B([1847]), .Y([1848]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11433 (.A([1848]), .Y([1849]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11434 (.A([1846]), .B([1849]), .Y([1850]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11435 (.A([1586]), .B([1850]), .X([1851]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11436 (.A([1851]), .Y([1852]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11437 (.A([1845]), .B([1852]), .Y([1853]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11438 (.A([1608]), .B([1839]), .X([1854]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11439 (.A([1607]), .B([1838]), .X([1855]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11440 (.A([1854]), .B([1855]), .Y([1856]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11441 (.A([1609]), .B([1856]), .Y([1857]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11442 (.A([1853]), .B([1854]), .X([1858]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11443 (.A([1853]), .B([1857]), .Y([1859]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11444 (.A([1858]), .B([1859]), .Y([1860]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11445 (.A([1558]), .B([1860]), .Y([1861]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11446 (.A([1844]), .B([1861]), .Y([1862]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11447 (.A([1843]), .B([1862]), .Y([1863]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11448 (.A([1842]), .B([1862]), .X([1864]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11449 (.A([1863]), .B([1864]), .Y([1865]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11450 (.A([1634]), .B([1640]), .Y([1866]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11451 (.A([1558]), .B([1866]), .Y([1867]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11452 (.A([1554]), .B([1867]), .X([1868]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11453 (.A([456]), .B([1867]), .Y([1869]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11454 (.A([1868]), .B([1869]), .Y([1870]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11455 (.A([1865]), .B([1870]), .X([1871]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11456 (.A([1863]), .B([1871]), .Y([1872]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11457 (.A([1813]), .B([1834]), .X([1873]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11458 (.A([1835]), .B([1873]), .Y([1874]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11459 (.A([1874]), .Y([1875]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11460 (.A([1872]), .B([1875]), .Y([1876]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11461 (.A([1835]), .B([1876]), .Y([1877]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11462 (.A([1783]), .B([1805]), .Y([1878]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11463 (.A([1806]), .B([1878]), .Y([1879]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11464 (.A([1879]), .Y([1880]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11465 (.A([1877]), .B([1880]), .Y([1881]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11466 (.A([1806]), .B([1881]), .Y([1882]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11467 (.A([1776]), .B([1882]), .Y([1883]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11468 (.A([1776]), .B([1882]), .X([1884]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11469 (.A([1883]), .B([1884]), .Y([1885]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11470 (.A([1886]), .B([1517]), .Y([1887]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11471 (.A([1887]), .Y([1888]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11472 (.A([1877]), .B([1880]), .X([1889]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11473 (.A([1881]), .B([1889]), .Y([1890]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11474 (.A([1872]), .B([1875]), .X([1891]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11475 (.A([1876]), .B([1891]), .Y([1892]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11476 (.A([1890]), .B([1892]), .Y([1893]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11477 (.A([1888]), .B([1893]), .Y([1894]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11478 (.A([1885]), .B([1894]), .X([1895]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11479 (.A([1773]), .B([1883]), .Y([1896]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11480 (.A([1896]), .Y([1897]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11481 (.A([1895]), .B([1897]), .Y([1898]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11482 (.A([1720]), .B([1743]), .X([1899]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11483 (.A([1744]), .B([1899]), .Y([1900]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11484 (.A([1900]), .Y([1901]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11485 (.A([1898]), .B([1901]), .Y([1902]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11486 (.A([1744]), .B([1902]), .Y([1903]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11487 (.A([1691]), .B([1712]), .Y([1904]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11488 (.A([1713]), .B([1904]), .Y([1905]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11489 (.A([1905]), .Y([1906]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11490 (.A([1903]), .B([1906]), .Y([1907]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11491 (.A([1713]), .B([1907]), .Y([1908]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11492 (.A([1661]), .B([1683]), .X([1909]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11493 (.A([1684]), .B([1909]), .Y([1910]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11494 (.A([1910]), .Y([1911]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11495 (.A([1908]), .B([1911]), .Y([1912]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11496 (.A([1684]), .B([1912]), .Y([1913]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11497 (.A([1631]), .B([1650]), .X([1914]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11498 (.A([1914]), .Y([1915]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11499 (.A([1646]), .B([1914]), .Y([1916]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11500 (.A([1913]), .B([1916]), .Y([1917]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11501 (.A([1913]), .B([1916]), .X([1918]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11502 (.A([1917]), .B([1918]), .Y([1919]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11503 (.A([433]), .B([1919]), .X([1920]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11504 (.A([1654]), .B([1920]), .Y([1921]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11505 (.A([1921]), .Y([1922]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11506 (.A([433]), .B([1923]), .Y([1924]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11507 (.A([39]), .B([1898]), .Y([1925]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11508 (.A([1924]), .B([1925]), .Y([1926]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11509 (.A([1865]), .B([1870]), .Y([1927]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11510 (.A([1871]), .B([1927]), .Y([1928]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11511 (.A([39]), .B([1928]), .Y([1929]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11512 (.A([39]), .B([516]), .X([1930]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11513 (.A([1929]), .B([1930]), .Y([1931]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11514 (.A([1931]), .Y([1932]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11515 (.A([39]), .B([286]), .X([1933]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11516 (.A([39]), .B([1892]), .Y([1934]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11517 (.A([1933]), .B([1934]), .Y([1935]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11518 (.A([1935]), .Y([1936]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11519 (.A([39]), .B([518]), .X([1937]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11520 (.A([39]), .B([1890]), .Y([1938]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11521 (.A([1937]), .B([1938]), .Y([1939]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11522 (.A([1939]), .Y([1940]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11523 (.A([39]), .B([145]), .X([1941]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11524 (.A([39]), .B([1885]), .Y([1942]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11525 (.A([1941]), .B([1942]), .Y([1943]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11526 (.A([1943]), .Y([1944]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11527 (.A([1898]), .B([1901]), .X([1945]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11528 (.A([1902]), .B([1945]), .Y([1946]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11529 (.A([39]), .B([1946]), .Y([1947]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11530 (.A([39]), .B([169]), .X([1948]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11531 (.A([1947]), .B([1948]), .Y([1949]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11532 (.A([1949]), .Y([1950]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11533 (.A([1903]), .B([1906]), .X([1951]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11534 (.A([1907]), .B([1951]), .Y([1952]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11535 (.A([39]), .B([191]), .X([1953]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11536 (.A([39]), .B([1952]), .Y([1954]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11537 (.A([1953]), .B([1954]), .Y([1955]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11538 (.A([1955]), .Y([1956]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11539 (.A([1908]), .B([1911]), .X([1957]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11540 (.A([1912]), .B([1957]), .Y([1958]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11541 (.A([39]), .B([213]), .X([1959]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11542 (.A([39]), .B([1958]), .Y([1960]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11543 (.A([1959]), .B([1960]), .Y([1961]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11544 (.A([1961]), .Y([1962]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11545 (.A([433]), .B([1963]), .Y([1964]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11546 (.A([39]), .B([1594]), .Y([1965]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11547 (.A([1964]), .B([1965]), .Y([1966]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11548 (.A([39]), .B([550]), .X([1967]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11549 (.A([1558]), .B([1853]), .X([1968]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11550 (.A([456]), .B([1556]), .Y([1969]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11551 (.A([1968]), .B([1969]), .Y([1970]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11552 (.A([1913]), .B([1915]), .X([1971]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11553 (.A([1646]), .B([1971]), .Y([1972]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11554 (.A([1970]), .B([1972]), .X([1973]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11555 (.A([1970]), .B([1972]), .Y([1974]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11556 (.A([1973]), .B([1974]), .Y([1975]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11557 (.A([1952]), .B([1958]), .Y([1976]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11558 (.A([1888]), .B([1976]), .Y([1977]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11559 (.A([39]), .B([1977]), .Y([1978]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11560 (.A([1920]), .B([1978]), .Y([1979]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11561 (.A([1975]), .B([1979]), .Y([1980]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11562 (.A([1967]), .B([1980]), .Y([1981]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11563 (.A([1981]), .Y([1982]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11564 (.A([1983]), .B([1125]), .X([1984]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11565 (.A([38]), .B([1985]), .Y([1986]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11566 (.A([1531]), .B([1986]), .X([1987]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11567 (.A([1988]), .B([1986]), .Y([1989]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11568 (.A([1987]), .B([1989]), .Y([1990]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11569 (.A([1984]), .B([1990]), .Y([1991]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11570 (.A([1991]), .Y([1992]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11571 (.A([456]), .B([1066]), .X([1993]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11572 (.A([1993]), .Y([1994]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11573 (.A([1995]), .B([1066]), .Y([1996]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11574 (.A([3]), .B([1996]), .Y([1997]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11575 (.A([1994]), .B([1997]), .X([1998]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11576 (.A([1404]), .B([1001]), .Y([1999]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11577 (.A([2000]), .B([1999]), .X([2001]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11578 (.A([696]), .B([1993]), .Y([2002]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11579 (.A([1531]), .B([695]), .Y([2003]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11580 (.A([2002]), .B([2003]), .Y([2004]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11581 (.A([1999]), .B([2004]), .Y([2005]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11582 (.A([2001]), .B([2005]), .Y([2006]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11583 (.A([1002]), .B([2006]), .X([2007]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11584 (.A([2007]), .Y([2008]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11585 (.A([2009]), .B([476]), .Y([2010]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11586 (.A([309]), .B([476]), .X([2011]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11587 (.A([2010]), .B([2011]), .Y([2012]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11588 (.A([660]), .B([2012]), .Y([2013]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11589 (.A([60]), .B([2014]), .Y([2015]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11590 (.A([2016]), .B([2009]), .Y([2017]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11591 (.A([2015]), .B([2017]), .Y([2018]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11592 (.A([2019]), .B([2018]), .Y([2020]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11593 (.A([2021]), .B([44]), .Y([2022]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11594 (.A([2020]), .B([2022]), .Y([2023]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11595 (.A([661]), .B([2023]), .Y([2024]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11596 (.A([2013]), .B([2024]), .Y([2025]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11597 (.A([469]), .B([2025]), .Y([2026]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11598 (.A([1015]), .B([469]), .X([2027]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11599 (.A([1125]), .B([2027]), .Y([2028]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11600 (.A([2028]), .Y([2029]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11601 (.A([2026]), .B([2029]), .Y([2030]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11602 (.A([1118]), .B([1183]), .X([2031]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11603 (.A([1193]), .B([2031]), .Y([2032]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11604 (.A([491]), .B([1601]), .X([2033]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11605 (.A([2033]), .Y([2034]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11606 (.A([456]), .B([2031]), .X([2035]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11607 (.A([2032]), .B([2035]), .Y([2036]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11608 (.A([2033]), .B([2036]), .X([116]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11609 (.A([602]), .B([2034]), .Y([2037]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11610 (.A([2038]), .B([2039]), .X([2040]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11611 (.A([150]), .B([2040]), .Y([2041]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11612 (.A([577]), .B([2041]), .Y([2042]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11613 (.A([2043]), .B([2039]), .X([2044]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11614 (.A([490]), .B([2044]), .Y([2045]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11615 (.A([516]), .B([2045]), .Y([2046]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11616 (.A([1274]), .B([1160]), .Y([2047]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11617 (.A([253]), .B([2047]), .Y([2048]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11618 (.A([675]), .B([1149]), .Y([2049]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11619 (.A([2042]), .B([2049]), .Y([2050]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11620 (.A([2046]), .B([2048]), .Y([2051]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11621 (.A([2051]), .Y([2052]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11622 (.A([2037]), .B([2052]), .Y([2053]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11623 (.A([2050]), .B([2053]), .X([108]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11624 (.A([718]), .B([2033]), .X([2054]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11625 (.A([286]), .B([2045]), .Y([2055]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11626 (.A([2055]), .Y([2056]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11627 (.A([531]), .B([2041]), .Y([2057]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11628 (.A([279]), .B([2047]), .Y([2058]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11629 (.A([721]), .B([1149]), .Y([2059]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11630 (.A([2058]), .B([2059]), .Y([2060]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11631 (.A([2060]), .Y([2061]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11632 (.A([2057]), .B([2061]), .Y([2062]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11633 (.A([2056]), .B([2062]), .X([2063]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11634 (.A([2063]), .Y([2064]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11635 (.A([2054]), .B([2064]), .Y([109]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11636 (.A([749]), .B([2033]), .X([2065]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11637 (.A([2009]), .B([2041]), .Y([2066]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11638 (.A([2066]), .Y([2067]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11639 (.A([518]), .B([2045]), .Y([2068]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11640 (.A([138]), .B([1149]), .Y([2069]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11641 (.A([303]), .B([2047]), .Y([2070]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11642 (.A([2069]), .B([2070]), .Y([2071]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11643 (.A([2071]), .Y([2072]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11644 (.A([2068]), .B([2072]), .Y([2073]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11645 (.A([2067]), .B([2073]), .X([2074]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11646 (.A([2074]), .Y([2075]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11647 (.A([2065]), .B([2075]), .Y([110]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11648 (.A([778]), .B([2033]), .X([2076]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11649 (.A([145]), .B([2045]), .Y([2077]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11650 (.A([474]), .B([2041]), .Y([2078]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11651 (.A([327]), .B([2047]), .Y([2079]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11652 (.A([142]), .B([1149]), .Y([2080]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11653 (.A([2078]), .B([2080]), .Y([2081]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11654 (.A([2077]), .B([2079]), .Y([2082]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11655 (.A([2082]), .Y([2083]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11656 (.A([2076]), .B([2083]), .Y([2084]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11657 (.A([2081]), .B([2084]), .X([111]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11658 (.A([807]), .B([2033]), .X([2085]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11659 (.A([169]), .B([2045]), .Y([2086]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11660 (.A([2086]), .Y([2087]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11661 (.A([349]), .B([2047]), .Y([2088]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11662 (.A([167]), .B([1149]), .Y([2089]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11663 (.A([2088]), .B([2089]), .Y([2090]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11664 (.A([1531]), .B([2040]), .X([2091]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11665 (.A([2092]), .B([150]), .X([2093]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11666 (.A([2091]), .B([2093]), .Y([2094]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11667 (.A([2090]), .B([2094]), .X([2095]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11668 (.A([2087]), .B([2095]), .X([2096]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11669 (.A([2096]), .Y([2097]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11670 (.A([2085]), .B([2097]), .Y([112]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11671 (.A([836]), .B([2033]), .X([2098]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11672 (.A([191]), .B([2045]), .Y([2099]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11673 (.A([2099]), .Y([2100]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11674 (.A([150]), .B([2091]), .Y([2101]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11675 (.A([189]), .B([1149]), .Y([2102]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11676 (.A([373]), .B([2047]), .Y([2103]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11677 (.A([2102]), .B([2103]), .Y([2104]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11678 (.A([2101]), .B([2104]), .X([2105]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11679 (.A([2100]), .B([2105]), .X([2106]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11680 (.A([2106]), .Y([2107]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11681 (.A([2098]), .B([2107]), .Y([113]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11682 (.A([865]), .B([2033]), .X([2108]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11683 (.A([213]), .B([2045]), .Y([2109]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11684 (.A([2110]), .B([2041]), .Y([2111]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11685 (.A([2111]), .Y([2112]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11686 (.A([211]), .B([1149]), .Y([2113]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11687 (.A([2113]), .Y([2114]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11688 (.A([396]), .B([2047]), .Y([2115]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11689 (.A([2109]), .B([2115]), .Y([2116]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11690 (.A([2114]), .B([2116]), .X([2117]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11691 (.A([2112]), .B([2117]), .X([2118]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11692 (.A([2118]), .Y([2119]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11693 (.A([2108]), .B([2119]), .Y([114]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11694 (.A([894]), .B([2033]), .X([2120]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11695 (.A([2121]), .B([2041]), .Y([2122]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11696 (.A([2122]), .Y([2123]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11697 (.A([236]), .B([2044]), .X([2124]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11698 (.A([499]), .B([2124]), .Y([2125]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11699 (.A([417]), .B([2047]), .Y([2126]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11700 (.A([232]), .B([1149]), .Y([2127]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11701 (.A([2126]), .B([2127]), .Y([2128]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11702 (.A([2125]), .B([2128]), .X([2129]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11703 (.A([2123]), .B([2129]), .X([2130]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11704 (.A([2130]), .Y([2131]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11705 (.A([2120]), .B([2131]), .Y([115]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11706 (.A([546]), .B([474]), .Y([2132]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11707 (.A([2132]), .Y([2133]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9277 (.A([2134]), .Y([705]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9278 (.A([2135]), .Y([595]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9279 (.A([2136]), .Y([587]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9280 (.A([2110]), .Y([1254]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9281 (.A([1988]), .Y([1983]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9282 (.A([60]), .Y([1531]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9283 (.A([462]), .Y([2137]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9284 (.A([2043]), .Y([2038]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9285 (.A([453]), .Y([459]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9286 (.A([2021]), .Y([2019]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9287 (.A([2014]), .Y([2016]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9288 (.A([2138]), .Y([2139]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9289 (.A([544]), .Y([484]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9290 (.A([39]), .Y([433]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9291 (.A([448]), .Y([1259]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9292 (.A([2121]), .Y([496]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9293 (.A([531]), .Y([1240]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9294 (.A([577]), .Y([1243]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9295 (.A([1006]), .Y([2140]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9296 (.A([1010]), .Y([2141]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9297 (.A([1013]), .Y([2142]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9298 (.A([1019]), .Y([2143]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9299 (.A([1023]), .Y([2144]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9300 (.A([1031]), .Y([2145]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9301 (.A([1036]), .Y([2146]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9302 (.A([2147]), .Y([1422]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9303 (.A([234]), .Y([236]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9304 (.A([516]), .Y([263]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9305 (.A([518]), .Y([309]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9306 (.A([169]), .Y([171]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9307 (.A([213]), .Y([215]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9308 (.A([44]), .Y([456]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9309 (.A([3]), .Y([1002]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9310 (.A([2148]), .Y([1247]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9311 (.A([1368]), .B([2149]), .X([488]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9312 (.A([488]), .Y([690]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9313 (.A([1216]), .B([2150]), .X([2151]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9314 (.A([1316]), .B([1346]), .X([608]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9315 (.A([2151]), .B([608]), .X([666]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9316 (.A([488]), .B([666]), .X([2039]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9317 (.A([1316]), .B([2152]), .X([2153]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9318 (.A([2151]), .B([2153]), .X([2154]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9319 (.A([1383]), .B([2155]), .X([614]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9320 (.A([614]), .Y([1123]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9321 (.A([2154]), .B([614]), .X([1274]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9322 (.A([1274]), .Y([2156]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9323 (.A([2039]), .B([1274]), .Y([1599]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9324 (.A([1368]), .B([1383]), .X([605]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9325 (.A([605]), .Y([2157]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9326 (.A([1216]), .B([1288]), .X([641]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9327 (.A([2153]), .B([641]), .X([1153]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9328 (.A([605]), .B([1153]), .X([1160]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9329 (.A([488]), .B([2154]), .X([1161]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9330 (.A([1288]), .B([2158]), .X([609]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9331 (.A([1346]), .B([2159]), .X([642]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9332 (.A([609]), .B([642]), .X([654]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9333 (.A([488]), .B([654]), .X([1132]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9334 (.A([1161]), .B([1132]), .Y([1264]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9335 (.A([2039]), .B([1160]), .Y([1563]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9336 (.A([2156]), .B([1264]), .X([2160]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9337 (.A([1563]), .B([2160]), .X([603]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9338 (.A([603]), .Y([719]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9339 (.A([2158]), .B([2150]), .X([2161]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9340 (.A([2153]), .B([2161]), .X([623]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9341 (.A([605]), .B([623]), .X([1125]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9342 (.A([2159]), .B([2152]), .X([2162]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9343 (.A([641]), .B([2162]), .X([2163]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9344 (.A([488]), .B([2163]), .X([629]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9345 (.A([1125]), .B([629]), .Y([2164]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9346 (.A([2161]), .B([2162]), .X([606]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9347 (.A([614]), .B([606]), .X([2165]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9348 (.A([2165]), .Y([697]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9349 (.A([488]), .B([1153]), .X([1188]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9350 (.A([2165]), .B([1188]), .Y([634]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9351 (.A([2151]), .B([2162]), .X([489]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9352 (.A([614]), .B([489]), .X([694]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9353 (.A([694]), .Y([1265]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9354 (.A([614]), .B([2163]), .X([1302]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9355 (.A([694]), .B([1302]), .Y([2166]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9356 (.A([2164]), .B([2166]), .X([2167]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9357 (.A([634]), .B([2167]), .X([2168]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9358 (.A([603]), .B([2168]), .X([2169]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9359 (.A([605]), .B([2163]), .X([1066]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9360 (.A([1066]), .Y([472]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9361 (.A([2169]), .B([472]), .X([2170]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9362 (.A([608]), .B([641]), .X([615]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9363 (.A([2155]), .B([2149]), .X([611]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9364 (.A([615]), .B([611]), .X([1133]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9365 (.A([608]), .B([2161]), .X([639]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9366 (.A([614]), .B([639]), .X([617]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9367 (.A([1133]), .B([617]), .Y([1359]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9368 (.A([605]), .B([489]), .X([1130]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9369 (.A([666]), .B([605]), .X([2171]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9370 (.A([1130]), .B([2171]), .Y([1276]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9371 (.A([1359]), .B([1276]), .X([1565]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9372 (.A([1565]), .Y([2172]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9373 (.A([1449]), .B([2172]), .Y([2173]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9374 (.A([2170]), .B([2173]), .X([2174]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9375 (.A([2175]), .B([1565]), .Y([2176]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9376 (.A([1410]), .B([472]), .Y([2177]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9377 (.A([2176]), .B([2177]), .Y([2178]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9378 (.A([2169]), .B([2178]), .X([2179]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9379 (.A([2179]), .Y([2180]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9380 (.A([2174]), .B([2180]), .Y([588]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9381 (.A([588]), .Y([737]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9382 (.A([1274]), .B([1302]), .Y([1335]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9383 (.A([1335]), .Y([1200]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9384 (.A([634]), .B([1335]), .X([1143]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9385 (.A([481]), .B([2181]), .Y([2182]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9386 (.A([1066]), .B([2182]), .X([2183]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9387 (.A([44]), .B([1066]), .Y([2184]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9388 (.A([2183]), .B([2184]), .Y([2185]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9389 (.A([1143]), .B([2185]), .X([2186]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9390 (.A([2164]), .B([2186]), .X([2187]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9391 (.A([39]), .B([2187]), .Y([2188]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9392 (.A([2188]), .Y([2189]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9393 (.A([1422]), .B([2170]), .X([2190]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9394 (.A([1386]), .B([472]), .Y([2191]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9395 (.A([2172]), .B([2191]), .Y([2192]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9396 (.A([2192]), .Y([2193]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9397 (.A([2190]), .B([2193]), .Y([600]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9398 (.A([600]), .Y([593]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9399 (.A([2189]), .B([600]), .Y([2194]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9400 (.A([737]), .B([2194]), .X([2195]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9401 (.A([2196]), .B([2197]), .X([2198]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9402 (.A([2199]), .B([2198]), .X([2200]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9403 (.A([1886]), .B([2196]), .X([2201]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9404 (.A([1923]), .B([2201]), .X([2202]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9405 (.A([2200]), .B([2202]), .Y([2203]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9406 (.A([1923]), .B([2197]), .X([2204]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9407 (.A([1886]), .B([2199]), .X([2205]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9408 (.A([2204]), .B([2205]), .Y([2206]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9409 (.A([2203]), .B([2206]), .X([2207]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9410 (.A([2196]), .B([2207]), .X([2208]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9411 (.A([44]), .B([2208]), .Y([2209]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9412 (.A([263]), .B([2209]), .Y([2210]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9413 (.A([263]), .B([2209]), .X([2211]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9414 (.A([2210]), .B([2211]), .Y([2212]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9415 (.A([1274]), .B([2212]), .Y([2213]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9416 (.A([39]), .B([2214]), .X([2215]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9417 (.A([433]), .B([20]), .X([2216]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9418 (.A([2215]), .B([2216]), .Y([567]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9419 (.A([567]), .Y([256]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9420 (.A([1274]), .B([256]), .X([2217]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9421 (.A([2217]), .Y([2218]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9422 (.A([2189]), .B([2213]), .Y([2219]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9423 (.A([2218]), .B([2219]), .X([2220]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9424 (.A([2195]), .B([2220]), .X([2221]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9425 (.A([597]), .B([2195]), .Y([2222]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9426 (.A([2221]), .B([2222]), .Y([2223]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9427 (.A([286]), .B([2203]), .Y([2224]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9428 (.A([286]), .B([2203]), .X([2225]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9429 (.A([2224]), .B([2225]), .Y([2226]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9430 (.A([2211]), .B([2226]), .Y([2227]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9431 (.A([2211]), .B([2226]), .X([2228]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9432 (.A([2227]), .B([2228]), .Y([2229]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9433 (.A([1274]), .B([2229]), .Y([2230]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9434 (.A([39]), .B([2231]), .X([2232]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9435 (.A([433]), .B([21]), .X([2233]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9436 (.A([2232]), .B([2233]), .Y([508]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9437 (.A([508]), .Y([281]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9438 (.A([1274]), .B([281]), .X([2234]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9439 (.A([2234]), .Y([2235]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9440 (.A([2189]), .B([2230]), .Y([2236]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9441 (.A([2235]), .B([2236]), .X([2237]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9442 (.A([2195]), .B([2237]), .X([2238]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9443 (.A([2134]), .B([2195]), .Y([2239]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9444 (.A([2238]), .B([2239]), .Y([2240]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9445 (.A([2224]), .B([2228]), .Y([2241]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9446 (.A([2241]), .Y([2242]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9447 (.A([309]), .B([2200]), .X([2243]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9448 (.A([309]), .B([2200]), .Y([2244]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9449 (.A([2243]), .B([2244]), .Y([2245]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9450 (.A([2242]), .B([2245]), .Y([2246]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9451 (.A([2242]), .B([2245]), .X([2247]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9452 (.A([2246]), .B([2247]), .Y([2248]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9453 (.A([1274]), .B([2248]), .Y([2249]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9454 (.A([39]), .B([2250]), .X([2251]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9455 (.A([433]), .B([22]), .X([2252]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9456 (.A([2251]), .B([2252]), .Y([1015]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9457 (.A([1015]), .Y([305]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9458 (.A([1274]), .B([305]), .X([2253]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9459 (.A([2189]), .B([2253]), .Y([2254]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9460 (.A([2254]), .Y([2255]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9461 (.A([2249]), .B([2255]), .Y([2256]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9462 (.A([2195]), .B([2256]), .X([2257]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9463 (.A([739]), .B([2195]), .Y([2258]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9464 (.A([2257]), .B([2258]), .Y([2259]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9465 (.A([2243]), .B([2247]), .Y([2260]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9466 (.A([145]), .B([2202]), .Y([2261]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9467 (.A([145]), .B([2202]), .X([2262]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9468 (.A([2261]), .B([2262]), .Y([2263]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9469 (.A([2263]), .Y([2264]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9470 (.A([2260]), .B([2264]), .Y([2265]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9471 (.A([2260]), .B([2264]), .X([2266]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9472 (.A([2265]), .B([2266]), .Y([2267]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9473 (.A([2156]), .B([2267]), .X([2268]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9474 (.A([39]), .B([2269]), .X([2270]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9475 (.A([433]), .B([23]), .X([2271]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9476 (.A([2270]), .B([2271]), .Y([468]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9477 (.A([468]), .Y([329]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9478 (.A([1274]), .B([329]), .X([2272]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9479 (.A([2189]), .B([2272]), .Y([2273]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9480 (.A([2273]), .Y([2274]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9481 (.A([2268]), .B([2274]), .Y([2275]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9482 (.A([2195]), .B([2275]), .X([2276]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9483 (.A([768]), .B([2195]), .Y([2277]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9484 (.A([2276]), .B([2277]), .Y([2278]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9485 (.A([2279]), .B([2198]), .X([2280]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9486 (.A([550]), .B([2201]), .X([2281]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9487 (.A([2280]), .B([2281]), .Y([2282]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9488 (.A([550]), .B([2197]), .X([2283]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9489 (.A([1886]), .B([2279]), .X([2284]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9490 (.A([2283]), .B([2284]), .Y([2285]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9491 (.A([2282]), .B([2285]), .X([2286]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9492 (.A([2196]), .B([2286]), .X([2287]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9493 (.A([44]), .B([2287]), .Y([2288]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9494 (.A([171]), .B([2288]), .Y([2289]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9495 (.A([171]), .B([2288]), .X([2290]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9496 (.A([2289]), .B([2290]), .Y([2291]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9497 (.A([1274]), .B([2291]), .Y([2292]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9498 (.A([39]), .B([24]), .Y([2293]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9499 (.A([433]), .B([2294]), .Y([2295]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9500 (.A([2293]), .B([2295]), .Y([352]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9501 (.A([1274]), .B([352]), .X([2296]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9502 (.A([2296]), .Y([2297]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9503 (.A([2189]), .B([2292]), .Y([2298]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9504 (.A([2297]), .B([2298]), .X([2299]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9505 (.A([2195]), .B([2299]), .X([2300]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9506 (.A([797]), .B([2195]), .Y([2301]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9507 (.A([2300]), .B([2301]), .Y([2302]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9508 (.A([191]), .B([2282]), .Y([2303]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9509 (.A([191]), .B([2282]), .X([2304]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9510 (.A([2303]), .B([2304]), .Y([2305]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9511 (.A([2290]), .B([2305]), .Y([2306]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9512 (.A([2290]), .B([2305]), .X([2307]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9513 (.A([2306]), .B([2307]), .Y([2308]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9514 (.A([1274]), .B([2308]), .Y([2309]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9515 (.A([39]), .B([2310]), .X([2311]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9516 (.A([433]), .B([25]), .X([2312]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9517 (.A([2311]), .B([2312]), .Y([1028]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9518 (.A([1028]), .Y([375]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9519 (.A([1274]), .B([375]), .X([2313]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9520 (.A([2313]), .Y([2314]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9521 (.A([2189]), .B([2309]), .Y([2315]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9522 (.A([2314]), .B([2315]), .X([2316]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9523 (.A([2195]), .B([2316]), .X([2317]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9524 (.A([826]), .B([2195]), .Y([2318]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9525 (.A([2317]), .B([2318]), .Y([2319]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9526 (.A([2303]), .B([2307]), .Y([2320]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9527 (.A([2320]), .Y([2321]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9528 (.A([215]), .B([2280]), .X([2322]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9529 (.A([215]), .B([2280]), .Y([2323]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9530 (.A([2322]), .B([2323]), .Y([2324]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9531 (.A([2321]), .B([2324]), .Y([2325]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9532 (.A([2321]), .B([2324]), .X([2326]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9533 (.A([2325]), .B([2326]), .Y([2327]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9534 (.A([1274]), .B([2327]), .Y([2328]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9535 (.A([39]), .B([2329]), .X([2330]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9536 (.A([433]), .B([26]), .X([2331]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9537 (.A([2330]), .B([2331]), .Y([1033]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9538 (.A([1033]), .Y([398]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9539 (.A([1274]), .B([398]), .X([2332]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9540 (.A([2189]), .B([2332]), .Y([2333]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9541 (.A([2333]), .Y([2334]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9542 (.A([2328]), .B([2334]), .Y([2335]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9543 (.A([2195]), .B([2335]), .X([2336]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9544 (.A([855]), .B([2195]), .Y([2337]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9545 (.A([2336]), .B([2337]), .Y([2338]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9546 (.A([2322]), .B([2326]), .Y([2339]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9547 (.A([234]), .B([2281]), .Y([2340]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9548 (.A([234]), .B([2281]), .X([2341]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9549 (.A([2340]), .B([2341]), .Y([2342]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9550 (.A([2339]), .B([2342]), .X([2343]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9551 (.A([2339]), .B([2342]), .Y([2344]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9552 (.A([2343]), .B([2344]), .Y([2345]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9553 (.A([1274]), .B([2345]), .Y([2346]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9554 (.A([433]), .B([2347]), .Y([2348]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9555 (.A([39]), .B([27]), .Y([585]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9556 (.A([2348]), .B([585]), .Y([419]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9557 (.A([1274]), .B([419]), .X([2349]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9558 (.A([2189]), .B([2349]), .Y([2350]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9559 (.A([2350]), .Y([2351]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9560 (.A([2346]), .B([2351]), .Y([2352]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9561 (.A([2195]), .B([2352]), .X([2353]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9562 (.A([884]), .B([2195]), .Y([2354]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9563 (.A([2353]), .B([2354]), .Y([2355]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9564 (.A([588]), .B([2194]), .X([2356]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9565 (.A([2135]), .B([2356]), .Y([2357]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9566 (.A([2220]), .B([2356]), .X([2358]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9567 (.A([2357]), .B([2358]), .Y([2359]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9568 (.A([707]), .B([2356]), .Y([2360]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9569 (.A([2237]), .B([2356]), .X([2361]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9570 (.A([2360]), .B([2361]), .Y([2362]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9571 (.A([736]), .B([2356]), .Y([2363]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9572 (.A([2256]), .B([2356]), .X([2364]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9573 (.A([2363]), .B([2364]), .Y([2365]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9574 (.A([2275]), .B([2356]), .X([2366]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9575 (.A([766]), .B([2356]), .Y([2367]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9576 (.A([2366]), .B([2367]), .Y([2368]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9577 (.A([2299]), .B([2356]), .X([2369]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9578 (.A([795]), .B([2356]), .Y([2370]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9579 (.A([2369]), .B([2370]), .Y([2371]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9580 (.A([2316]), .B([2356]), .X([2372]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9581 (.A([824]), .B([2356]), .Y([2373]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9582 (.A([2372]), .B([2373]), .Y([2374]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9583 (.A([2335]), .B([2356]), .X([2375]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9584 (.A([853]), .B([2356]), .Y([2376]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9585 (.A([2375]), .B([2376]), .Y([2377]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9586 (.A([882]), .B([2356]), .Y([2378]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9587 (.A([2352]), .B([2356]), .X([2379]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9588 (.A([2378]), .B([2379]), .Y([2380]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9589 (.A([588]), .B([593]), .Y([482]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9590 (.A([2188]), .B([482]), .X([2381]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9591 (.A([590]), .B([2381]), .Y([2382]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9592 (.A([2220]), .B([2381]), .X([2383]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9593 (.A([2382]), .B([2383]), .Y([2384]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9594 (.A([2237]), .B([2381]), .X([2385]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9595 (.A([711]), .B([2381]), .Y([2386]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9596 (.A([2385]), .B([2386]), .Y([2387]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9597 (.A([743]), .B([2381]), .Y([2388]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9598 (.A([2256]), .B([2381]), .X([2389]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9599 (.A([2388]), .B([2389]), .Y([2390]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9600 (.A([2275]), .B([2381]), .X([2391]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9601 (.A([775]), .B([2381]), .Y([2392]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9602 (.A([2391]), .B([2392]), .Y([2393]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9603 (.A([801]), .B([2381]), .Y([2394]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9604 (.A([2299]), .B([2381]), .X([2395]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9605 (.A([2394]), .B([2395]), .Y([2396]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9606 (.A([2316]), .B([2381]), .X([2397]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9607 (.A([830]), .B([2381]), .Y([2398]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9608 (.A([2397]), .B([2398]), .Y([2399]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9609 (.A([2335]), .B([2381]), .X([2400]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9610 (.A([859]), .B([2381]), .Y([2401]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9611 (.A([2400]), .B([2401]), .Y([2402]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9612 (.A([2352]), .B([2381]), .X([2403]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9613 (.A([891]), .B([2381]), .Y([2404]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9614 (.A([2403]), .B([2404]), .Y([2405]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9615 (.A([588]), .B([600]), .X([715]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9616 (.A([2188]), .B([715]), .X([2406]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9617 (.A([2136]), .B([2406]), .Y([2407]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9618 (.A([2220]), .B([2406]), .X([2408]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9619 (.A([2407]), .B([2408]), .Y([2409]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9620 (.A([2237]), .B([2406]), .X([2410]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9621 (.A([714]), .B([2406]), .Y([2411]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9622 (.A([2410]), .B([2411]), .Y([2412]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9623 (.A([2256]), .B([2406]), .X([2413]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9624 (.A([746]), .B([2406]), .Y([2414]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9625 (.A([2413]), .B([2414]), .Y([2415]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9626 (.A([772]), .B([2406]), .Y([2416]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9627 (.A([2275]), .B([2406]), .X([2417]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9628 (.A([2416]), .B([2417]), .Y([2418]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9629 (.A([2299]), .B([2406]), .X([2419]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9630 (.A([804]), .B([2406]), .Y([2420]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9631 (.A([2419]), .B([2420]), .Y([2421]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9632 (.A([2316]), .B([2406]), .X([2422]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9633 (.A([833]), .B([2406]), .Y([2423]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9634 (.A([2422]), .B([2423]), .Y([2424]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9635 (.A([2335]), .B([2406]), .X([2425]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9636 (.A([862]), .B([2406]), .Y([2426]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9637 (.A([2425]), .B([2426]), .Y([2427]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9638 (.A([888]), .B([2406]), .Y([2428]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9639 (.A([2352]), .B([2406]), .X([2429]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9640 (.A([2428]), .B([2429]), .Y([2430]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9641 (.A([1963]), .B([550]), .X([2431]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9642 (.A([1963]), .B([550]), .Y([2432]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9643 (.A([2431]), .B([2432]), .Y([2433]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9644 (.A([1513]), .B([234]), .Y([2434]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9645 (.A([1513]), .B([234]), .X([2435]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9646 (.A([2434]), .B([2435]), .Y([2436]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9647 (.A([2433]), .B([2436]), .Y([2437]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9648 (.A([2433]), .B([2436]), .X([2438]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9649 (.A([2437]), .B([2438]), .Y([2439]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9650 (.A([2139]), .B([546]), .Y([2440]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9651 (.A([2440]), .Y([2441]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9652 (.A([2439]), .B([2441]), .Y([2442]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9653 (.A([2138]), .B([456]), .Y([2443]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9654 (.A([2137]), .B([2443]), .Y([2444]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9655 (.A([2444]), .Y([2445]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9656 (.A([2442]), .B([2445]), .Y([2446]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9657 (.A([2446]), .Y([2447]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9658 (.A([462]), .B([213]), .Y([2448]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9659 (.A([642]), .B([2161]), .X([2449]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9660 (.A([488]), .B([2449]), .X([469]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9661 (.A([469]), .Y([542]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9662 (.A([472]), .B([469]), .Y([2450]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9663 (.A([2450]), .Y([466]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9664 (.A([2448]), .B([466]), .Y([2451]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9665 (.A([2447]), .B([2451]), .X([2452]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9666 (.A([609]), .B([2162]), .X([2453]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9667 (.A([605]), .B([2453]), .X([1113]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9668 (.A([1113]), .Y([1517]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9669 (.A([511]), .B([1517]), .Y([2454]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9670 (.A([472]), .B([2454]), .X([494]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9671 (.A([469]), .B([494]), .Y([2455]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9672 (.A([2455]), .Y([501]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9673 (.A([2137]), .B([1066]), .X([476]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9674 (.A([2138]), .B([546]), .X([2456]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9675 (.A([462]), .B([2456]), .X([2457]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9676 (.A([472]), .B([2457]), .Y([2458]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9677 (.A([1254]), .B([2458]), .Y([2459]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9678 (.A([501]), .B([2459]), .Y([2460]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9679 (.A([398]), .B([2455]), .Y([2461]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9680 (.A([2460]), .B([2461]), .Y([2462]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9681 (.A([2452]), .B([2462]), .Y([2463]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9682 (.A([2463]), .Y([2464]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9683 (.A([433]), .B([1066]), .X([1404]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9684 (.A([1404]), .Y([1387]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9685 (.A([462]), .B([1404]), .Y([2465]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9686 (.A([2000]), .B([398]), .X([2466]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9687 (.A([37]), .B([2467]), .Y([2468]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9688 (.A([1988]), .B([37]), .X([2092]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9689 (.A([1988]), .B([2467]), .X([2469]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9690 (.A([2092]), .B([2469]), .Y([2470]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9691 (.A([1983]), .B([2468]), .Y([2471]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9692 (.A([2000]), .B([2145]), .Y([2472]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9693 (.A([2466]), .B([2472]), .Y([2473]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9694 (.A([2471]), .B([2473]), .X([2474]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9695 (.A([2474]), .Y([2475]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9696 (.A([2000]), .B([419]), .X([2476]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9697 (.A([2000]), .B([2146]), .Y([2477]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9698 (.A([2470]), .B([2477]), .Y([2478]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9699 (.A([2478]), .Y([2479]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9700 (.A([2476]), .B([2479]), .Y([1455]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9701 (.A([1455]), .Y([2480]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9702 (.A([2000]), .B([352]), .X([2481]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9703 (.A([2000]), .B([2144]), .Y([2482]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9704 (.A([2481]), .B([2482]), .Y([2483]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9705 (.A([2471]), .B([2483]), .X([1349]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9706 (.A([1349]), .Y([1174]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9707 (.A([44]), .B([2471]), .Y([2484]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9708 (.A([1349]), .B([2484]), .Y([1094]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9709 (.A([1094]), .Y([1058]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9710 (.A([1455]), .B([2484]), .Y([450]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9711 (.A([450]), .Y([1497]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9712 (.A([1349]), .B([1497]), .Y([1087]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9713 (.A([1087]), .Y([1083]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9714 (.A([2000]), .B([1028]), .X([2485]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9715 (.A([2000]), .B([1026]), .Y([2486]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9716 (.A([2485]), .B([2486]), .Y([2487]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9717 (.A([2470]), .B([2487]), .Y([1506]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9718 (.A([1094]), .B([1506]), .X([1049]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9719 (.A([1087]), .B([1506]), .X([1046]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9720 (.A([2474]), .B([2484]), .Y([445]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9721 (.A([1046]), .B([445]), .X([1040]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9722 (.A([2000]), .B([281]), .X([2488]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9723 (.A([2000]), .B([2141]), .Y([2489]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9724 (.A([2470]), .B([2489]), .Y([2490]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9725 (.A([2490]), .Y([2491]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9726 (.A([2488]), .B([2491]), .Y([2492]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9727 (.A([2492]), .Y([2493]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9728 (.A([2000]), .B([256]), .X([2494]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9729 (.A([2000]), .B([2140]), .Y([2495]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9730 (.A([2494]), .B([2495]), .Y([2496]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9731 (.A([2471]), .B([2496]), .X([2497]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9732 (.A([2497]), .Y([1097]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9733 (.A([2484]), .B([2497]), .Y([2498]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9734 (.A([2493]), .B([2498]), .X([1055]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9735 (.A([1055]), .Y([1431]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9736 (.A([2000]), .B([329]), .X([2499]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9737 (.A([2000]), .B([2143]), .Y([2500]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9738 (.A([2499]), .B([2500]), .Y([2501]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9739 (.A([2471]), .B([2501]), .X([2502]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9740 (.A([2000]), .B([305]), .X([2503]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9741 (.A([2000]), .B([2142]), .Y([2504]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9742 (.A([2470]), .B([2504]), .Y([2505]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9743 (.A([2505]), .Y([2506]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9744 (.A([2503]), .B([2506]), .Y([1061]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9745 (.A([2484]), .B([1061]), .Y([1069]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9746 (.A([2502]), .B([1069]), .X([1395]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9747 (.A([1055]), .B([1395]), .X([1047]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9748 (.A([1404]), .B([1047]), .X([2507]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9749 (.A([1040]), .B([2507]), .X([2508]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9750 (.A([2465]), .B([2508]), .Y([2509]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9751 (.A([2043]), .B([1404]), .Y([2510]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9752 (.A([1083]), .B([1506]), .Y([1076]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9753 (.A([2475]), .B([1076]), .X([1101]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9754 (.A([2507]), .B([1101]), .X([2511]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9755 (.A([2510]), .B([2511]), .Y([2512]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9756 (.A([554]), .B([1404]), .Y([2513]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9757 (.A([2474]), .B([1497]), .Y([1460]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9758 (.A([2484]), .B([1506]), .Y([440]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9759 (.A([440]), .Y([2514]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9760 (.A([1349]), .B([440]), .X([1412]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9761 (.A([2507]), .B([1412]), .X([2515]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9762 (.A([1460]), .B([2515]), .X([2516]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9763 (.A([2513]), .B([2516]), .Y([2517]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9764 (.A([552]), .B([1404]), .Y([2518]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9765 (.A([1094]), .B([440]), .Y([2519]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9766 (.A([2507]), .B([2519]), .X([2520]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9767 (.A([1460]), .B([2520]), .X([2521]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9768 (.A([2518]), .B([2521]), .Y([2522]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9769 (.A([453]), .B([1404]), .Y([2523]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9770 (.A([450]), .B([445]), .Y([1477]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9771 (.A([2515]), .B([1477]), .X([2524]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9772 (.A([2523]), .B([2524]), .Y([2525]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9773 (.A([454]), .B([1404]), .Y([2526]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9774 (.A([2520]), .B([1477]), .X([2527]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9775 (.A([2526]), .B([2527]), .Y([2528]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9776 (.A([2021]), .B([1404]), .Y([2529]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9777 (.A([2474]), .B([450]), .X([1050]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9778 (.A([2515]), .B([1050]), .X([2530]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9779 (.A([2529]), .B([2530]), .Y([2531]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9780 (.A([2014]), .B([1404]), .Y([2532]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9781 (.A([2520]), .B([1050]), .X([2533]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9782 (.A([2532]), .B([2533]), .Y([2534]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9783 (.A([2138]), .B([1404]), .Y([2535]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9784 (.A([1455]), .B([445]), .X([1413]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9785 (.A([1413]), .Y([2536]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9786 (.A([2520]), .B([1413]), .X([2537]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9787 (.A([2535]), .B([2537]), .Y([2538]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9788 (.A([511]), .B([1404]), .Y([2539]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9789 (.A([2498]), .B([1061]), .X([2540]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9790 (.A([1055]), .B([1061]), .X([2541]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9791 (.A([1040]), .B([2541]), .X([1463]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9792 (.A([1404]), .B([1463]), .X([2542]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9793 (.A([2539]), .B([2542]), .Y([2543]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9794 (.A([1523]), .B([1404]), .Y([2544]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9795 (.A([2492]), .B([2498]), .X([1072]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9796 (.A([1395]), .B([1072]), .X([1085]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9797 (.A([1061]), .B([1072]), .X([2545]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9798 (.A([1085]), .B([2545]), .Y([2546]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9799 (.A([1404]), .B([450]), .X([2547]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9800 (.A([2547]), .Y([2548]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9801 (.A([2546]), .B([2548]), .Y([2549]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9802 (.A([2514]), .B([2549]), .X([2550]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9803 (.A([450]), .B([1085]), .X([2551]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9804 (.A([2544]), .B([2550]), .Y([2552]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9805 (.A([1050]), .B([1072]), .X([1464]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9806 (.A([1404]), .B([1464]), .X([2553]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9807 (.A([1555]), .B([1404]), .Y([2554]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9808 (.A([2553]), .B([2554]), .Y([2555]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9809 (.A([2484]), .B([2502]), .Y([1062]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9810 (.A([1062]), .Y([2556]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9811 (.A([2541]), .B([2556]), .X([1052]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9812 (.A([1052]), .Y([1043]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9813 (.A([1455]), .B([1094]), .X([1041]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9814 (.A([2474]), .B([1041]), .X([2557]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9815 (.A([1052]), .B([2557]), .X([2558]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9816 (.A([1055]), .B([1477]), .X([1393]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9817 (.A([1174]), .B([1062]), .X([2559]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9818 (.A([1393]), .B([2559]), .X([2560]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9819 (.A([2558]), .B([2560]), .Y([1484]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9820 (.A([2492]), .B([1097]), .Y([1073]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9821 (.A([2475]), .B([1506]), .Y([1088]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9822 (.A([1073]), .B([1088]), .X([1495]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9823 (.A([1497]), .B([1495]), .X([2561]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9824 (.A([1387]), .B([2561]), .Y([2562]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9825 (.A([1484]), .B([2562]), .X([2563]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9826 (.A([484]), .B([1404]), .Y([2564]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9827 (.A([2563]), .B([2564]), .Y([2565]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9828 (.A([2565]), .Y([2566]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9829 (.A([539]), .B([1404]), .Y([2567]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9830 (.A([2549]), .B([2567]), .Y([2568]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9831 (.A([1160]), .B([1066]), .Y([2569]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9832 (.A([39]), .B([2569]), .Y([2570]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9833 (.A([546]), .B([2570]), .Y([2571]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9834 (.A([445]), .B([440]), .Y([1456]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9835 (.A([1073]), .B([2570]), .X([2572]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9836 (.A([1456]), .B([2572]), .X([2573]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9837 (.A([2571]), .B([2573]), .Y([2574]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9838 (.A([1886]), .B([2570]), .Y([2575]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9839 (.A([474]), .B([1497]), .Y([2576]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9840 (.A([2573]), .B([2576]), .X([2577]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9841 (.A([2575]), .B([2577]), .Y([2578]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9842 (.A([1477]), .B([2545]), .X([1473]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9843 (.A([2514]), .B([1473]), .X([2579]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9844 (.A([1047]), .B([2557]), .X([2580]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9845 (.A([2579]), .B([2580]), .Y([2581]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9846 (.A([1387]), .B([2581]), .Y([2582]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9847 (.A([1543]), .B([1404]), .Y([2583]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9848 (.A([2582]), .B([2583]), .Y([2584]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9849 (.A([1506]), .B([1413]), .X([1397]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9850 (.A([1404]), .B([1397]), .X([2585]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9851 (.A([1525]), .B([1404]), .Y([2586]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9852 (.A([2585]), .B([2586]), .Y([2587]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9853 (.A([1196]), .B([1404]), .Y([2588]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9854 (.A([1387]), .B([1413]), .Y([2589]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9855 (.A([2545]), .B([2589]), .X([2590]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9856 (.A([2588]), .B([2590]), .Y([2591]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9857 (.A([2540]), .B([1073]), .Y([2592]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9858 (.A([1193]), .B([1404]), .Y([2593]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9859 (.A([2536]), .B([2592]), .Y([2594]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9860 (.A([1404]), .B([440]), .X([2595]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9861 (.A([2594]), .B([2595]), .X([2596]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9862 (.A([2593]), .B([2596]), .Y([2597]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9863 (.A([1061]), .B([2556]), .Y([1056]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9864 (.A([1073]), .B([1056]), .X([1064]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9865 (.A([1058]), .B([1064]), .X([1219]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9866 (.A([1395]), .B([1073]), .X([1095]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9867 (.A([1387]), .B([1095]), .Y([2598]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9868 (.A([1413]), .B([1072]), .X([2599]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9869 (.A([2599]), .Y([1438]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9870 (.A([1349]), .B([1413]), .X([2600]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9871 (.A([2545]), .B([2600]), .X([2601]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9872 (.A([1219]), .B([2601]), .Y([2602]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9873 (.A([2598]), .B([2602]), .X([2603]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9874 (.A([2175]), .B([1387]), .X([2604]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9875 (.A([2603]), .B([2604]), .Y([2605]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9876 (.A([2605]), .Y([2606]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9877 (.A([481]), .B([1387]), .X([2607]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9878 (.A([1047]), .B([2551]), .Y([2608]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9879 (.A([1058]), .B([2608]), .Y([2609]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9880 (.A([2609]), .Y([2610]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9881 (.A([2540]), .B([1085]), .Y([2611]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9882 (.A([1349]), .B([1397]), .X([1445]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9883 (.A([1097]), .B([1413]), .X([2612]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9884 (.A([2502]), .B([440]), .X([1436]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9885 (.A([1069]), .B([1436]), .X([2613]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9886 (.A([2480]), .B([1506]), .Y([2614]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9887 (.A([2614]), .Y([2615]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9888 (.A([1094]), .B([2614]), .X([1389]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9889 (.A([1041]), .B([1088]), .X([1428]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9890 (.A([1085]), .B([1428]), .X([1479]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9891 (.A([1479]), .Y([1406]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9892 (.A([1073]), .B([2615]), .X([2616]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9893 (.A([1445]), .B([1479]), .Y([2617]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9894 (.A([2611]), .B([2617]), .Y([2618]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9895 (.A([1413]), .B([2613]), .X([2619]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9896 (.A([2498]), .B([2619]), .X([2620]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9897 (.A([2616]), .B([2620]), .Y([2621]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9898 (.A([2621]), .Y([2622]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9899 (.A([2618]), .B([2622]), .Y([2623]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9900 (.A([1049]), .B([2612]), .X([2624]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9901 (.A([1387]), .B([2624]), .Y([2625]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9902 (.A([2623]), .B([2625]), .X([2626]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9903 (.A([2610]), .B([2626]), .X([2627]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9904 (.A([2607]), .B([2627]), .Y([2628]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9905 (.A([2628]), .Y([2629]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9906 (.A([1066]), .B([2471]), .X([2630]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9907 (.A([2151]), .B([642]), .X([621]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9908 (.A([605]), .B([621]), .X([172]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9909 (.A([172]), .Y([148]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9910 (.A([583]), .B([550]), .X([2631]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9911 (.A([583]), .B([550]), .Y([2632]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9912 (.A([2631]), .B([2632]), .Y([1184]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9913 (.A([148]), .B([1184]), .Y([1331]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9914 (.A([2630]), .B([1331]), .Y([2633]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9915 (.A([1125]), .B([1113]), .Y([2634]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9916 (.A([605]), .B([2449]), .X([264]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9917 (.A([264]), .Y([287]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9918 (.A([488]), .B([2453]), .X([2635]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9919 (.A([264]), .B([2635]), .Y([2636]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9920 (.A([2634]), .B([2636]), .X([2637]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9921 (.A([2633]), .B([2637]), .X([2638]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9922 (.A([44]), .B([172]), .Y([1578]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9923 (.A([472]), .B([1578]), .X([2639]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9924 (.A([2639]), .Y([2640]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9925 (.A([614]), .B([2449]), .X([2641]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9926 (.A([2153]), .B([609]), .X([631]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9927 (.A([488]), .B([631]), .X([2642]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9928 (.A([2641]), .B([2642]), .Y([1115]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9929 (.A([614]), .B([631]), .X([1126]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9930 (.A([1126]), .Y([2643]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9931 (.A([1115]), .B([2643]), .X([650]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9932 (.A([605]), .B([654]), .X([1295]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9933 (.A([1295]), .Y([1262]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9934 (.A([666]), .B([615]), .Y([691]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9935 (.A([2157]), .B([691]), .Y([1201]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9936 (.A([1295]), .B([1201]), .Y([1144]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9937 (.A([650]), .B([1144]), .X([2644]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9938 (.A([2640]), .B([2644]), .X([2645]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9939 (.A([2638]), .B([2645]), .X([2646]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9940 (.A([614]), .B([2453]), .X([2647]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9941 (.A([2635]), .B([2647]), .Y([1119]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9942 (.A([650]), .B([1119]), .X([146]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9943 (.A([2154]), .B([605]), .X([150]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9944 (.A([150]), .Y([199]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9945 (.A([1066]), .B([172]), .Y([2648]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9946 (.A([199]), .B([2648]), .X([1141]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9947 (.A([287]), .B([1141]), .X([2649]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9948 (.A([146]), .B([2649]), .X([2650]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9949 (.A([2630]), .B([2650]), .Y([254]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9950 (.A([287]), .B([254]), .X([143]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9951 (.A([675]), .B([143]), .Y([2651]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9952 (.A([516]), .B([146]), .Y([2652]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9953 (.A([1066]), .B([2470]), .X([2653]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9954 (.A([2653]), .Y([153]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9955 (.A([678]), .B([153]), .Y([2654]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9956 (.A([263]), .B([172]), .X([681]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9957 (.A([2654]), .B([681]), .Y([2655]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9958 (.A([2655]), .Y([2656]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9959 (.A([2652]), .B([2656]), .Y([2657]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9960 (.A([2657]), .Y([2658]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9961 (.A([2651]), .B([2658]), .Y([2659]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9962 (.A([2646]), .B([2659]), .Y([2660]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9963 (.A([2660]), .Y([2661]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9964 (.A([2646]), .B([2659]), .X([2662]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9965 (.A([2660]), .B([2662]), .Y([2663]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9966 (.A([39]), .B([2663]), .Y([2664]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9967 (.A([675]), .B([39]), .X([2665]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9968 (.A([2664]), .B([2665]), .Y([2666]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9969 (.A([2666]), .Y([2667]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9970 (.A([721]), .B([143]), .Y([2668]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9971 (.A([286]), .B([146]), .Y([2669]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9972 (.A([724]), .B([153]), .Y([2670]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9973 (.A([286]), .B([148]), .Y([2671]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9974 (.A([2671]), .Y([729]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9975 (.A([2672]), .B([199]), .Y([2673]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9976 (.A([2670]), .B([2673]), .Y([2674]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9977 (.A([2669]), .B([2671]), .Y([2675]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9978 (.A([2674]), .B([2675]), .X([2676]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9979 (.A([2676]), .Y([2677]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9980 (.A([2668]), .B([2677]), .Y([2678]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9981 (.A([2661]), .B([2678]), .Y([2679]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9982 (.A([2679]), .Y([132]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9983 (.A([2661]), .B([2678]), .X([2680]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9984 (.A([2679]), .B([2680]), .Y([2681]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9985 (.A([39]), .B([2681]), .Y([2682]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9986 (.A([39]), .B([721]), .X([2683]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9987 (.A([2682]), .B([2683]), .Y([2684]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9988 (.A([2684]), .Y([2685]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9989 (.A([138]), .B([143]), .Y([130]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9990 (.A([518]), .B([146]), .Y([2686]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9991 (.A([2686]), .Y([127]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9992 (.A([753]), .B([153]), .Y([2687]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9993 (.A([309]), .B([172]), .X([2688]));
  sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9994 (.A([2688]), .Y([124]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9995 (.A([1531]), .B([1995]), .Y([2689]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9996 (.A([1995]), .B([2690]), .X([2691]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9997 (.A([2689]), .B([2691]), .Y([2692]));
  sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9998 (.A([150]), .B([2692]), .X([2693]));
  sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9999 (.A([2687]), .B([2693]), .Y([125]));
  sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:40:hilomap_worker$12031 (.HI([2694]));
  sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:40:hilomap_worker$8815 (.HI([60]));
  sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:48:hilomap_worker$8817 (.LO([44]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11708 (.A([531]), .Y([2695]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11709 (.A([577]), .Y([2696]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11710 (.A([2110]), .Y([2697]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11711 (.A([2121]), .Y([2698]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11712 (.A([44]), .Y([2699]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11713 (.A([60]), .Y([2700]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11714 (.A([60]), .Y([2701]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11715 (.A([44]), .Y([2702]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11716 (.A([60]), .Y([2703]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11717 (.A([44]), .Y([2704]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11718 (.A([60]), .Y([2705]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11719 (.A([60]), .Y([2706]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11720 (.A([44]), .Y([2707]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11721 (.A([60]), .Y([2708]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11722 (.A([44]), .Y([2709]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11723 (.A([44]), .Y([2710]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11724 (.A([44]), .Y([2711]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11725 (.A([60]), .Y([2712]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11726 (.A([44]), .Y([2713]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11727 (.A([60]), .Y([2714]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11728 (.A([44]), .Y([2715]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11729 (.A([44]), .Y([2716]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11730 (.A([60]), .Y([2717]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11731 (.A([44]), .Y([2718]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11732 (.A([44]), .Y([2719]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11733 (.A([60]), .Y([2720]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11734 (.A([44]), .Y([2721]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11735 (.A([44]), .Y([2722]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11736 (.A([60]), .Y([2723]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11737 (.A([44]), .Y([2724]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11738 (.A([44]), .Y([2725]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11739 (.A([60]), .Y([2726]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11740 (.A([60]), .Y([2727]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11741 (.A([44]), .Y([2728]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11742 (.A([44]), .Y([2729]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11743 (.A([44]), .Y([2730]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11744 (.A([60]), .Y([2731]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11745 (.A([60]), .Y([2732]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11746 (.A([44]), .Y([2733]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11747 (.A([44]), .Y([2734]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11748 (.A([60]), .Y([2735]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11749 (.A([60]), .Y([2736]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11750 (.A([60]), .Y([2737]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11751 (.A([44]), .Y([2738]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11752 (.A([60]), .Y([2739]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11753 (.A([44]), .Y([2740]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11754 (.A([2741]), .Y([2742]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11755 (.A([60]), .Y([2743]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11756 (.A([44]), .Y([2744]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11757 (.A([44]), .Y([2745]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11758 (.A([44]), .Y([2746]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11759 (.A([60]), .Y([2747]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11760 (.A([44]), .Y([2748]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11761 (.A([44]), .Y([2749]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11762 (.A([60]), .Y([2750]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11763 (.A([44]), .Y([2751]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11764 (.A([60]), .Y([2752]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11765 (.A([60]), .Y([2753]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11766 (.A([44]), .Y([2754]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11767 (.A([44]), .Y([2755]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11768 (.A([60]), .Y([2756]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11769 (.A([44]), .Y([2757]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11770 (.A([60]), .Y([2758]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11771 (.A([60]), .Y([2759]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11772 (.A([44]), .Y([2760]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11773 (.A([60]), .Y([2761]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11774 (.A([44]), .Y([2762]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11775 (.A([44]), .Y([2763]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11776 (.A([60]), .Y([2764]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11777 (.A([60]), .Y([2765]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11778 (.A([44]), .Y([2766]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11779 (.A([60]), .Y([2767]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11780 (.A([60]), .Y([2768]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11781 (.A([60]), .Y([2769]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11782 (.A([44]), .Y([2770]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11783 (.A([60]), .Y([2771]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11784 (.A([44]), .Y([2772]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11785 (.A([60]), .Y([2773]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11786 (.A([60]), .Y([2774]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11787 (.A([44]), .Y([2775]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11788 (.A([44]), .Y([2776]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11789 (.A([60]), .Y([2777]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11790 (.A([44]), .Y([2778]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11791 (.A([60]), .Y([2779]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11792 (.A([44]), .Y([2780]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11793 (.A([44]), .Y([2781]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11794 (.A([44]), .Y([2782]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11795 (.A([60]), .Y([2783]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11796 (.A([44]), .Y([2784]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11797 (.A([60]), .Y([2785]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11798 (.A([60]), .Y([2786]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11799 (.A([60]), .Y([2787]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11800 (.A([60]), .Y([2788]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11801 (.A([44]), .Y([2789]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11802 (.A([44]), .Y([2790]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11803 (.A([60]), .Y([2791]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11804 (.A([44]), .Y([2792]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11805 (.A([60]), .Y([2793]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11806 (.A([60]), .Y([2794]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11807 (.A([44]), .Y([2795]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11808 (.A([44]), .Y([2796]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11809 (.A([60]), .Y([2797]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11810 (.A([60]), .Y([2798]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11811 (.A([44]), .Y([2799]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11812 (.A([60]), .Y([2800]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11813 (.A([60]), .Y([2801]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11814 (.A([60]), .Y([2802]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11815 (.A([44]), .Y([2803]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11816 (.A([44]), .Y([2804]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11817 (.A([44]), .Y([2805]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11818 (.A([60]), .Y([2806]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11819 (.A([60]), .Y([2807]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11820 (.A([60]), .Y([2808]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11821 (.A([44]), .Y([2809]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11822 (.A([60]), .Y([2810]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11823 (.A([60]), .Y([2811]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11824 (.A([44]), .Y([2812]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11825 (.A([60]), .Y([2813]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11826 (.A([60]), .Y([2814]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11827 (.A([44]), .Y([2815]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11828 (.A([44]), .Y([2816]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11829 (.A([44]), .Y([2817]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11830 (.A([44]), .Y([2818]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11831 (.A([44]), .Y([2819]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11832 (.A([44]), .Y([2820]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11833 (.A([60]), .Y([2821]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11834 (.A([60]), .Y([2822]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11835 (.A([60]), .Y([2823]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11836 (.A([60]), .Y([2824]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11837 (.A([60]), .Y([2825]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11838 (.A([60]), .Y([2826]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11839 (.A([44]), .Y([2827]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11840 (.A([44]), .Y([2828]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11841 (.A([60]), .Y([2829]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11842 (.A([44]), .Y([2830]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11843 (.A([44]), .Y([2831]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11844 (.A([44]), .Y([2832]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11845 (.A([60]), .Y([2833]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11846 (.A([44]), .Y([2834]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11847 (.A([60]), .Y([2835]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11848 (.A([60]), .Y([2836]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11849 (.A([60]), .Y([2837]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11850 (.A([44]), .Y([2838]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11851 (.A([60]), .Y([2839]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11852 (.A([60]), .Y([2840]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11853 (.A([44]), .Y([2841]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11854 (.A([60]), .Y([2842]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11855 (.A([44]), .Y([2843]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11856 (.A([44]), .Y([2844]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11857 (.A([44]), .Y([2845]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11858 (.A([60]), .Y([2846]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11859 (.A([44]), .Y([2847]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11860 (.A([60]), .Y([2848]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11861 (.A([44]), .Y([2849]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11862 (.A([60]), .Y([2850]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11863 (.A([60]), .Y([2851]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11864 (.A([44]), .Y([2852]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11865 (.A([44]), .Y([2853]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11866 (.A([60]), .Y([2854]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11867 (.A([44]), .Y([2855]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11868 (.A([60]), .Y([2856]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11869 (.A([44]), .Y([2857]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11870 (.A([44]), .Y([2858]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11871 (.A([44]), .Y([2859]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11872 (.A([60]), .Y([2860]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11873 (.A([44]), .Y([2861]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11874 (.A([44]), .Y([2862]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11875 (.A([44]), .Y([2863]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11876 (.A([44]), .Y([2864]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11877 (.A([44]), .Y([2865]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11878 (.A([60]), .Y([2866]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11879 (.A([44]), .Y([2867]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11880 (.A([60]), .Y([2868]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11881 (.A([60]), .Y([2869]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11882 (.A([60]), .Y([2870]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11883 (.A([60]), .Y([2871]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11884 (.A([44]), .Y([2872]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11885 (.A([44]), .Y([2873]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11886 (.A([60]), .Y([2874]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11887 (.A([1196]), .Y([2875]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11888 (.A([562]), .Y([2876]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11889 (.A([44]), .Y([2877]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11890 (.A([1196]), .Y([2878]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11891 (.A([2879]), .Y([2880]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11892 (.A([44]), .Y([2881]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11893 (.A([60]), .Y([2882]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11894 (.A([44]), .Y([2883]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11895 (.A([44]), .Y([2884]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11896 (.A([60]), .Y([2885]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11897 (.A([60]), .Y([2886]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11898 (.A([44]), .Y([2887]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11899 (.A([44]), .Y([2888]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11900 (.A([44]), .Y([2889]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11901 (.A([44]), .Y([2890]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11902 (.A([60]), .Y([2891]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11903 (.A([44]), .Y([2892]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11904 (.A([44]), .Y([2893]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11905 (.A([44]), .Y([2894]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11906 (.A([44]), .Y([2895]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11907 (.A([44]), .Y([2896]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11908 (.A([60]), .Y([2897]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11909 (.A([44]), .Y([2898]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11910 (.A([44]), .Y([2899]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11911 (.A([44]), .Y([2900]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11912 (.A([60]), .Y([2901]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11913 (.A([60]), .Y([2902]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11914 (.A([44]), .Y([2903]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11915 (.A([60]), .Y([2904]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11916 (.A([60]), .Y([2905]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11917 (.A([60]), .Y([2906]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11918 (.A([60]), .Y([2907]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11919 (.A([60]), .Y([2908]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11920 (.A([60]), .Y([2909]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11921 (.A([60]), .Y([2910]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11922 (.A([60]), .Y([2911]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11923 (.A([60]), .Y([2912]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11924 (.A([60]), .Y([2913]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11925 (.A([60]), .Y([2914]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11926 (.A([60]), .Y([2915]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11927 (.A([60]), .Y([2916]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11928 (.A([675]), .Y([2917]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11929 (.A([721]), .Y([2918]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11930 (.A([138]), .Y([2919]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11931 (.A([142]), .Y([2920]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11932 (.A([167]), .Y([2921]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11933 (.A([189]), .Y([2922]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11934 (.A([211]), .Y([2923]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11935 (.A([232]), .Y([2924]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11936 (.A([516]), .Y([2925]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11937 (.A([286]), .Y([2926]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11938 (.A([518]), .Y([2927]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11939 (.A([145]), .Y([2928]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11940 (.A([169]), .Y([2929]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11941 (.A([191]), .Y([2930]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11942 (.A([213]), .Y([2931]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11943 (.A([234]), .Y([2932]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11944 (.A([516]), .Y([2933]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11945 (.A([286]), .Y([2934]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11946 (.A([518]), .Y([2935]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11947 (.A([145]), .Y([2936]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11948 (.A([169]), .Y([2937]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11949 (.A([191]), .Y([2938]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11950 (.A([213]), .Y([2939]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11951 (.A([234]), .Y([2940]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11952 (.A([258]), .Y([2941]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11953 (.A([283]), .Y([2942]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11954 (.A([307]), .Y([2943]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11955 (.A([331]), .Y([2944]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11956 (.A([355]), .Y([2945]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11957 (.A([378]), .Y([2946]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11958 (.A([400]), .Y([2947]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11959 (.A([421]), .Y([2948]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11960 (.A([516]), .Y([2949]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11961 (.A([286]), .Y([2950]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11962 (.A([518]), .Y([2951]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11963 (.A([145]), .Y([2952]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11964 (.A([169]), .Y([2953]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11965 (.A([191]), .Y([2954]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11966 (.A([213]), .Y([2955]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11967 (.A([234]), .Y([2956]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11968 (.A([256]), .Y([2957]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11969 (.A([281]), .Y([2958]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11970 (.A([305]), .Y([2959]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11971 (.A([329]), .Y([2960]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11972 (.A([352]), .Y([2961]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11973 (.A([375]), .Y([2962]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11974 (.A([398]), .Y([2963]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11975 (.A([419]), .Y([2964]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11976 (.A([234]), .Y([2965]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11977 (.A([44]), .Y([45]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11978 (.A([44]), .Y([54]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11979 (.A([44]), .Y([55]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11980 (.A([44]), .Y([56]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11981 (.A([44]), .Y([57]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11982 (.A([44]), .Y([58]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11983 (.A([44]), .Y([59]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11984 (.A([60]), .Y([61]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11985 (.A([60]), .Y([62]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11986 (.A([60]), .Y([63]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11987 (.A([44]), .Y([46]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11988 (.A([60]), .Y([64]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11989 (.A([60]), .Y([65]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11990 (.A([60]), .Y([66]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11991 (.A([60]), .Y([67]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11992 (.A([44]), .Y([68]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11993 (.A([44]), .Y([69]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11994 (.A([44]), .Y([70]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11995 (.A([44]), .Y([71]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11996 (.A([44]), .Y([72]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11997 (.A([44]), .Y([73]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11998 (.A([44]), .Y([47]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11999 (.A([44]), .Y([74]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12000 (.A([44]), .Y([75]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12001 (.A([44]), .Y([76]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12002 (.A([60]), .Y([77]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12003 (.A([60]), .Y([78]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12004 (.A([60]), .Y([79]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12005 (.A([60]), .Y([80]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12006 (.A([60]), .Y([81]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12007 (.A([60]), .Y([82]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12008 (.A([60]), .Y([83]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12009 (.A([44]), .Y([48]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12010 (.A([44]), .Y([49]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12011 (.A([44]), .Y([50]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12012 (.A([44]), .Y([51]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12013 (.A([44]), .Y([52]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12014 (.A([44]), .Y([53]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12015 (.A([44]), .Y([100]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12016 (.A([44]), .Y([101]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12017 (.A([44]), .Y([102]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12018 (.A([44]), .Y([103]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12019 (.A([44]), .Y([104]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12020 (.A([44]), .Y([105]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12021 (.A([44]), .Y([106]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12022 (.A([44]), .Y([107]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12023 (.A([44]), .Y([117]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12024 (.A([44]), .Y([118]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12025 (.A([44]), .Y([119]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12026 (.A([44]), .Y([120]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12027 (.A([44]), .Y([121]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12028 (.A([44]), .Y([122]));
  sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12029 (.A([44]), .Y([123]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4105 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2223]), .Q([597]), .Q_N([2966]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4106 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2240]), .Q([2134]), .Q_N([2967]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4107 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2259]), .Q([739]), .Q_N([2968]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4108 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2278]), .Q([768]), .Q_N([2969]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4109 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2302]), .Q([797]), .Q_N([2970]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4110 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2319]), .Q([826]), .Q_N([2971]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4111 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2338]), .Q([855]), .Q_N([2972]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4112 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2355]), .Q([884]), .Q_N([2973]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4907 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2359]), .Q([2135]), .Q_N([2974]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4908 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2362]), .Q([707]), .Q_N([2975]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4909 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2365]), .Q([736]), .Q_N([2976]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4910 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2368]), .Q([766]), .Q_N([2977]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4911 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2371]), .Q([795]), .Q_N([2978]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4912 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2374]), .Q([824]), .Q_N([2979]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4913 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2377]), .Q([853]), .Q_N([2980]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4914 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2380]), .Q([882]), .Q_N([2981]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4931 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2384]), .Q([590]), .Q_N([2982]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4932 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2387]), .Q([711]), .Q_N([2983]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4933 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2390]), .Q([743]), .Q_N([2984]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4934 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2393]), .Q([775]), .Q_N([2985]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4935 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2396]), .Q([801]), .Q_N([2986]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4936 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2399]), .Q([830]), .Q_N([2987]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4937 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2402]), .Q([859]), .Q_N([2988]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4938 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2405]), .Q([891]), .Q_N([2989]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4979 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2409]), .Q([2136]), .Q_N([2990]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4980 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2412]), .Q([714]), .Q_N([2991]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4981 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2415]), .Q([746]), .Q_N([2992]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4982 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2418]), .Q([772]), .Q_N([2993]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4983 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2421]), .Q([804]), .Q_N([2994]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4984 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2424]), .Q([833]), .Q_N([2995]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4985 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2427]), .Q([862]), .Q_N([2996]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4986 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2430]), .Q([888]), .Q_N([2997]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5134 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2464]), .Q([2110]), .Q_N([1251]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5135 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1992]), .Q([1988]), .Q_N([2690]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5136 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([38]), .Q([2998]), .Q_N([1985]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5137 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2509]), .Q([462]), .Q_N([2181]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5138 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2512]), .Q([2043]), .Q_N([2999]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5139 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2517]), .Q([554]), .Q_N([3000]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5140 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2522]), .Q([552]), .Q_N([3001]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5141 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2525]), .Q([453]), .Q_N([3002]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5142 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2528]), .Q([454]), .Q_N([3003]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5143 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2531]), .Q([2021]), .Q_N([3004]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5144 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2534]), .Q([2014]), .Q_N([3005]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5145 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2538]), .Q([2138]), .Q_N([3006]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5146 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2543]), .Q([511]), .Q_N([3007]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5151 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2552]), .Q([1523]), .Q_N([3008]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5152 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2555]), .Q([1555]), .Q_N([3009]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5153 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2566]), .Q([544]), .Q_N([3010]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5154 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2568]), .Q([539]), .Q_N([3011]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5155 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2574]), .Q([546]), .Q_N([3012]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5156 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2578]), .Q([1886]), .Q_N([2197]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5157 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2584]), .Q([1543]), .Q_N([3013]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5158 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2587]), .Q([1525]), .Q_N([3014]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5159 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2591]), .Q([1196]), .Q_N([562]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5160 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2597]), .Q([1193]), .Q_N([3015]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5161 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2606]), .Q([2175]), .Q_N([3016]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5166 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2629]), .Q([481]), .Q_N([3017]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5167 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2667]), .Q([675]), .Q_N([3018]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5168 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2685]), .Q([721]), .Q_N([3019]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5169 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([141]), .Q([138]), .Q_N([3020]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5170 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([166]), .Q([142]), .Q_N([3021]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5171 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([188]), .Q([167]), .Q_N([3022]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5172 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([210]), .Q([189]), .Q_N([3023]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5173 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([231]), .Q([211]), .Q_N([3024]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5174 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([252]), .Q([232]), .Q_N([3025]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5175 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([278]), .Q([253]), .Q_N([3026]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5176 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([302]), .Q([279]), .Q_N([3027]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5177 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([326]), .Q([303]), .Q_N([3028]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5178 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([348]), .Q([327]), .Q_N([3029]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5179 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([372]), .Q([349]), .Q_N([3030]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5180 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([395]), .Q([373]), .Q_N([3031]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5181 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([416]), .Q([396]), .Q_N([3032]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5182 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([437]), .Q([417]), .Q_N([3033]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5183 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1998]), .Q([1995]), .Q_N([2672]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5189 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([256]), .Q([2214]), .Q_N([3034]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5190 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([281]), .Q([2231]), .Q_N([3035]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5191 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([305]), .Q([2250]), .Q_N([3036]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5192 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([329]), .Q([2269]), .Q_N([3037]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5193 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([352]), .Q([2294]), .Q_N([3038]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5194 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([375]), .Q([2310]), .Q_N([3039]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5195 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([398]), .Q([2329]), .Q_N([3040]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5196 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([419]), .Q([2347]), .Q_N([3041]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5197 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([442]), .Q([438]), .Q_N([1238]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5198 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([447]), .Q([443]), .Q_N([1232]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5199 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([452]), .Q([448]), .Q_N([2148]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5200 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2008]), .Q([2000]), .Q_N([3042]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5201 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([480]), .Q([474]), .Q_N([3043]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5202 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([507]), .Q([2121]), .Q_N([1249]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5203 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2030]), .Q([2009]), .Q_N([2467]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5204 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([538]), .Q([531]), .Q_N([1235]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5205 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([582]), .Q([577]), .Q_N([1230]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5206 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([586]), .Q([583]), .Q_N([3044]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5207 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([704]), .Q([678]), .Q_N([3045]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5208 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([735]), .Q([724]), .Q_N([3046]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5209 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([765]), .Q([753]), .Q_N([3047]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5210 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([794]), .Q([152]), .Q_N([3048]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5211 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([823]), .Q([175]), .Q_N([3049]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5212 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([852]), .Q([194]), .Q_N([3050]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5213 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([881]), .Q([218]), .Q_N([3051]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5214 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([908]), .Q([239]), .Q_N([3052]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5215 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([2133]), .Q([3053]), .Q_N([2196]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5216 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([921]), .Q([258]), .Q_N([3054]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5217 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([932]), .Q([283]), .Q_N([3055]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5218 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([943]), .Q([307]), .Q_N([3056]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5219 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([954]), .Q([331]), .Q_N([3057]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5220 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([965]), .Q([355]), .Q_N([3058]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5221 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([976]), .Q([378]), .Q_N([3059]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5222 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([989]), .Q([400]), .Q_N([3060]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5223 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1000]), .Q([421]), .Q_N([3061]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5224 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1008]), .Q([1006]), .Q_N([3062]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5225 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1012]), .Q([1010]), .Q_N([3063]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5226 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1017]), .Q([1013]), .Q_N([3064]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5227 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1021]), .Q([1019]), .Q_N([3065]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5228 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1025]), .Q([1023]), .Q_N([3066]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5229 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1030]), .Q([1026]), .Q_N([3067]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5230 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1035]), .Q([1031]), .Q_N([3068]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5231 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1039]), .Q([1036]), .Q_N([3069]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5232 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1218]), .Q([1216]), .Q_N([2158]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5233 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1291]), .Q([1288]), .Q_N([2150]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5234 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1318]), .Q([1316]), .Q_N([2159]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5235 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1348]), .Q([1346]), .Q_N([2152]), .RESET_B([2694]), .SET_B([3]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5236 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1370]), .Q([1368]), .Q_N([2155]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5237 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1385]), .Q([1383]), .Q_N([2149]), .RESET_B([3]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8804 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1409]), .Q([1386]), .Q_N([3070]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8805 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1421]), .Q([1410]), .Q_N([3071]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8806 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1444]), .Q([2147]), .Q_N([3072]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8807 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1452]), .Q([1449]), .Q_N([3073]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8808 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1472]), .Q([1453]), .Q_N([3074]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8809 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1490]), .Q([1488]), .Q_N([3075]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8810 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1503]), .Q([1491]), .Q_N([3076]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8811 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1512]), .Q([1504]), .Q_N([3077]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7456 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1653]), .Q([1513]), .Q_N([3078]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7679 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1922]), .Q([234]), .Q_N([3079]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7680 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1926]), .Q([1923]), .Q_N([2199]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7681 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1932]), .Q([516]), .Q_N([3080]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7682 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1936]), .Q([286]), .Q_N([3081]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7683 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1940]), .Q([518]), .Q_N([3082]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7684 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1944]), .Q([145]), .Q_N([3083]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7685 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1950]), .Q([169]), .Q_N([3084]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7686 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1956]), .Q([191]), .Q_N([3085]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7687 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1962]), .Q([213]), .Q_N([3086]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7689 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1966]), .Q([1963]), .Q_N([3087]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7690 (.CLK(clk_buf_T35Y0__R3_BUF_0_out), .D([1982]), .Q([550]), .Q_N([2279]), .RESET_B([2694]), .SET_B([2694]));
  sky130_fd_sc_hd__clkbuf_4 T0Y0__R0_BUF_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R0_INV_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y0__R1_BUF_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R1_INV_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R2_INV_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y0__R2_INV_1 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y0__R3_BUF_0 (.A(tie_lo_T0Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y10__R0_BUF_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R0_INV_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y10__R1_BUF_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R1_INV_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R2_INV_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y10__R2_INV_1 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y10__R3_BUF_0 (.A(tie_lo_T0Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y11__R0_BUF_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R0_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y11__R1_BUF_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R1_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R2_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y11__R2_INV_1 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y11__R3_BUF_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y12__R0_BUF_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R0_INV_0 (.A(tie_lo_T0Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y12__R1_BUF_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R1_INV_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R2_INV_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y12__R2_INV_1 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y12__R3_BUF_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y13__R0_BUF_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R0_INV_0 (.A(tie_lo_T0Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y13__R1_BUF_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R1_INV_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R2_INV_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y13__R2_INV_1 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y13__R3_BUF_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y14__R0_BUF_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R0_INV_0 (.A(tie_lo_T0Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y14__R1_BUF_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R1_INV_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R2_INV_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y14__R2_INV_1 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y14__R3_BUF_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y15__R0_BUF_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R0_INV_0 (.A(tie_lo_T0Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y15__R1_BUF_0 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R1_INV_0 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R2_INV_0 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y15__R2_INV_1 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y15__R3_BUF_0 (.A(tie_lo_T0Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y16__R0_BUF_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R0_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y16__R1_BUF_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R1_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R2_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y16__R2_INV_1 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y16__R3_BUF_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y17__R0_BUF_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R0_INV_0 (.A(tie_lo_T0Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y17__R1_BUF_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R1_INV_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R2_INV_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y17__R2_INV_1 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y17__R3_BUF_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y18__R0_BUF_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R0_INV_0 (.A(tie_lo_T0Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y18__R1_BUF_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R1_INV_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R2_INV_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y18__R2_INV_1 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y18__R3_BUF_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y19__R0_BUF_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R0_INV_0 (.A(tie_lo_T0Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y19__R1_BUF_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R1_INV_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R2_INV_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y19__R2_INV_1 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y19__R3_BUF_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y1__R0_BUF_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R0_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y1__R1_BUF_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R1_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R2_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y1__R2_INV_1 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y1__R3_BUF_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y20__R0_BUF_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R0_INV_0 (.A(tie_lo_T0Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y20__R1_BUF_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R1_INV_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R2_INV_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y20__R2_INV_1 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y20__R3_BUF_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y21__R0_BUF_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R0_INV_0 (.A(tie_lo_T0Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y21__R1_BUF_0 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R1_INV_0 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R2_INV_0 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y21__R2_INV_1 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y21__R3_BUF_0 (.A(tie_lo_T0Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y22__R0_BUF_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R0_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y22__R1_BUF_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R1_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R2_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y22__R2_INV_1 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y22__R3_BUF_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y23__R0_BUF_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R0_INV_0 (.A(tie_lo_T0Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y23__R1_BUF_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R1_INV_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R2_INV_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y23__R2_INV_1 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y23__R3_BUF_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y24__R0_BUF_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R0_INV_0 (.A(tie_lo_T0Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y24__R1_BUF_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R1_INV_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R2_INV_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y24__R2_INV_1 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y24__R3_BUF_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y25__R0_BUF_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R0_INV_0 (.A(tie_lo_T0Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y25__R1_BUF_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R1_INV_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R2_INV_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y25__R2_INV_1 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y25__R3_BUF_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y26__R0_BUF_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R0_INV_0 (.A(tie_lo_T0Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y26__R1_BUF_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R1_INV_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R2_INV_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y26__R2_INV_1 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y26__R3_BUF_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y27__R0_BUF_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R0_INV_0 (.A(tie_lo_T0Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y27__R1_BUF_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R1_INV_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R2_INV_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y27__R2_INV_1 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y27__R3_BUF_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y28__R0_BUF_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R0_INV_0 (.A(tie_lo_T0Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y28__R1_BUF_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R1_INV_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R2_INV_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y28__R2_INV_1 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y28__R3_BUF_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y29__R0_BUF_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R0_INV_0 (.A(tie_lo_T0Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y29__R1_BUF_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R1_INV_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R2_INV_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y29__R2_INV_1 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y29__R3_BUF_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y2__R0_BUF_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R0_INV_0 (.A(tie_lo_T0Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y2__R1_BUF_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R1_INV_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R2_INV_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y2__R2_INV_1 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y2__R3_BUF_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y30__R0_BUF_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R0_INV_0 (.A(tie_lo_T0Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y30__R1_BUF_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R1_INV_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R2_INV_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y30__R2_INV_1 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y30__R3_BUF_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y31__R0_BUF_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R0_INV_0 (.A(tie_lo_T0Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y31__R1_BUF_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R1_INV_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R2_INV_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y31__R2_INV_1 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y31__R3_BUF_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y32__R0_BUF_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R0_INV_0 (.A(tie_lo_T0Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y32__R1_BUF_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R1_INV_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R2_INV_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y32__R2_INV_1 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y32__R3_BUF_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y33__R0_BUF_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R0_INV_0 (.A(tie_lo_T0Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y33__R1_BUF_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R1_INV_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R2_INV_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y33__R2_INV_1 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y33__R3_BUF_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y34__R0_BUF_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R0_INV_0 (.A(tie_lo_T0Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y34__R1_BUF_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R1_INV_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R2_INV_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y34__R2_INV_1 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y34__R3_BUF_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y35__R0_BUF_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R0_INV_0 (.A(tie_lo_T0Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y35__R1_BUF_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R1_INV_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R2_INV_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y35__R2_INV_1 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y35__R3_BUF_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y36__R0_BUF_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R0_INV_0 (.A(tie_lo_T0Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y36__R1_BUF_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R1_INV_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R2_INV_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y36__R2_INV_1 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y36__R3_BUF_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y37__R0_BUF_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R0_INV_0 (.A(tie_lo_T0Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y37__R1_BUF_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R1_INV_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R2_INV_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y37__R2_INV_1 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y37__R3_BUF_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y38__R0_BUF_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R0_INV_0 (.A(tie_lo_T0Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y38__R1_BUF_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R1_INV_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R2_INV_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y38__R2_INV_1 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y38__R3_BUF_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y39__R0_BUF_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R0_INV_0 (.A(tie_lo_T0Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y39__R1_BUF_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R1_INV_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R2_INV_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y39__R2_INV_1 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y39__R3_BUF_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y3__R0_BUF_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R0_INV_0 (.A(tie_lo_T0Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y3__R1_BUF_0 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R1_INV_0 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R2_INV_0 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y3__R2_INV_1 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y3__R3_BUF_0 (.A(tie_lo_T0Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y40__R0_BUF_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R0_INV_0 (.A(tie_lo_T0Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y40__R1_BUF_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R1_INV_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R2_INV_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y40__R2_INV_1 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y40__R3_BUF_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y41__R0_BUF_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R0_INV_0 (.A(tie_lo_T0Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y41__R1_BUF_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R1_INV_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R2_INV_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y41__R2_INV_1 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y41__R3_BUF_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y42__R0_BUF_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R0_INV_0 (.A(tie_lo_T0Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y42__R1_BUF_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R1_INV_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R2_INV_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y42__R2_INV_1 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y42__R3_BUF_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y43__R0_BUF_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R0_INV_0 (.A(tie_lo_T0Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y43__R1_BUF_0 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R1_INV_0 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R2_INV_0 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y43__R2_INV_1 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y43__R3_BUF_0 (.A(tie_lo_T0Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y44__R0_BUF_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R0_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y44__R1_BUF_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R1_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R2_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y44__R2_INV_1 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y44__R3_BUF_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y45__R0_BUF_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R0_INV_0 (.A(tie_lo_T0Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y45__R1_BUF_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R1_INV_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R2_INV_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y45__R2_INV_1 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y45__R3_BUF_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y46__R0_BUF_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R0_INV_0 (.A(tie_lo_T0Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y46__R1_BUF_0 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R1_INV_0 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R2_INV_0 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y46__R2_INV_1 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y46__R3_BUF_0 (.A(tie_lo_T0Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y47__R0_BUF_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R0_INV_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y47__R1_BUF_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R1_INV_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R2_INV_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y47__R2_INV_1 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y47__R3_BUF_0 (.A(tie_lo_T0Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y48__R0_BUF_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R0_INV_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y48__R1_BUF_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R1_INV_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R2_INV_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y48__R2_INV_1 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y48__R3_BUF_0 (.A(tie_lo_T0Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y49__R0_BUF_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R0_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y49__R1_BUF_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R1_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R2_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y49__R2_INV_1 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y49__R3_BUF_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y4__R0_BUF_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R0_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y4__R1_BUF_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R1_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R2_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y4__R2_INV_1 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y4__R3_BUF_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y50__R0_BUF_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R0_INV_0 (.A(tie_lo_T0Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y50__R1_BUF_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R1_INV_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R2_INV_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y50__R2_INV_1 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y50__R3_BUF_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y51__R0_BUF_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R0_INV_0 (.A(tie_lo_T0Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y51__R1_BUF_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R1_INV_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R2_INV_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y51__R2_INV_1 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y51__R3_BUF_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y52__R0_BUF_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R0_INV_0 (.A(tie_lo_T0Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y52__R1_BUF_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R1_INV_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R2_INV_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y52__R2_INV_1 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y52__R3_BUF_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y53__R0_BUF_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R0_INV_0 (.A(tie_lo_T0Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y53__R1_BUF_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R1_INV_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R2_INV_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y53__R2_INV_1 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y53__R3_BUF_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y54__R0_BUF_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R0_INV_0 (.A(tie_lo_T0Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y54__R1_BUF_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R1_INV_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R2_INV_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y54__R2_INV_1 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y54__R3_BUF_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y55__R0_BUF_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R0_INV_0 (.A(tie_lo_T0Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y55__R1_BUF_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R1_INV_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R2_INV_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y55__R2_INV_1 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y55__R3_BUF_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y56__R0_BUF_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R0_INV_0 (.A(tie_lo_T0Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y56__R1_BUF_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R1_INV_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R2_INV_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y56__R2_INV_1 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y56__R3_BUF_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y57__R0_BUF_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R0_INV_0 (.A(tie_lo_T0Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y57__R1_BUF_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R1_INV_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R2_INV_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y57__R2_INV_1 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y57__R3_BUF_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y58__R0_BUF_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R0_INV_0 (.A(tie_lo_T0Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y58__R1_BUF_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R1_INV_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R2_INV_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y58__R2_INV_1 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y58__R3_BUF_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y59__R0_BUF_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R0_INV_0 (.A(tie_lo_T0Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y59__R1_BUF_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R1_INV_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R2_INV_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y59__R2_INV_1 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y59__R3_BUF_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y5__R0_BUF_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R0_INV_0 (.A(tie_lo_T0Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y5__R1_BUF_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R1_INV_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R2_INV_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y5__R2_INV_1 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y5__R3_BUF_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y60__R0_BUF_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R0_INV_0 (.A(tie_lo_T0Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y60__R1_BUF_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R1_INV_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R2_INV_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y60__R2_INV_1 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y60__R3_BUF_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y61__R0_BUF_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R0_INV_0 (.A(tie_lo_T0Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y61__R1_BUF_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R1_INV_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R2_INV_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y61__R2_INV_1 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y61__R3_BUF_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y62__R0_BUF_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R0_INV_0 (.A(tie_lo_T0Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y62__R1_BUF_0 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R1_INV_0 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R2_INV_0 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y62__R2_INV_1 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y62__R3_BUF_0 (.A(tie_lo_T0Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y63__R0_BUF_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R0_INV_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y63__R1_BUF_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R1_INV_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R2_INV_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y63__R2_INV_1 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y63__R3_BUF_0 (.A(tie_lo_T0Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y64__R0_BUF_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R0_INV_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y64__R1_BUF_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R1_INV_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R2_INV_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y64__R2_INV_1 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y64__R3_BUF_0 (.A(tie_lo_T0Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y65__R0_BUF_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R0_INV_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y65__R1_BUF_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R1_INV_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R2_INV_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y65__R2_INV_1 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y65__R3_BUF_0 (.A(tie_lo_T0Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y66__R0_BUF_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R0_INV_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y66__R1_BUF_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R1_INV_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R2_INV_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y66__R2_INV_1 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y66__R3_BUF_0 (.A(tie_lo_T0Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y67__R0_BUF_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R0_INV_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y67__R1_BUF_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R1_INV_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R2_INV_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y67__R2_INV_1 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y67__R3_BUF_0 (.A(tie_lo_T0Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y68__R0_BUF_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R0_INV_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y68__R1_BUF_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R1_INV_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R2_INV_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y68__R2_INV_1 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y68__R3_BUF_0 (.A(tie_lo_T0Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y69__R0_BUF_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R0_INV_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y69__R1_BUF_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R1_INV_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R2_INV_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y69__R2_INV_1 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y69__R3_BUF_0 (.A(tie_lo_T0Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y6__R0_BUF_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R0_INV_0 (.A(tie_lo_T0Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y6__R1_BUF_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R1_INV_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R2_INV_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y6__R2_INV_1 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y6__R3_BUF_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y70__R0_BUF_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R0_INV_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y70__R1_BUF_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R1_INV_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R2_INV_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y70__R2_INV_1 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y70__R3_BUF_0 (.A(tie_lo_T0Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y71__R0_BUF_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R0_INV_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y71__R1_BUF_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R1_INV_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R2_INV_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y71__R2_INV_1 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y71__R3_BUF_0 (.A(tie_lo_T0Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y72__R0_BUF_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R0_INV_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y72__R1_BUF_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R1_INV_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R2_INV_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y72__R2_INV_1 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y72__R3_BUF_0 (.A(tie_lo_T0Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y73__R0_BUF_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R0_INV_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y73__R1_BUF_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R1_INV_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R2_INV_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y73__R2_INV_1 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y73__R3_BUF_0 (.A(tie_lo_T0Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y74__R0_BUF_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R0_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y74__R1_BUF_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R1_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R2_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y74__R2_INV_1 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y74__R3_BUF_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y75__R0_BUF_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R0_INV_0 (.A(tie_lo_T0Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y75__R1_BUF_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R1_INV_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R2_INV_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y75__R2_INV_1 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y75__R3_BUF_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y76__R0_BUF_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R0_INV_0 (.A(tie_lo_T0Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y76__R1_BUF_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R1_INV_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R2_INV_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y76__R2_INV_1 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y76__R3_BUF_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y77__R0_BUF_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R0_INV_0 (.A(tie_lo_T0Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y77__R1_BUF_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R1_INV_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R2_INV_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y77__R2_INV_1 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y77__R3_BUF_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y78__R0_BUF_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R0_INV_0 (.A(tie_lo_T0Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y78__R1_BUF_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R1_INV_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R2_INV_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y78__R2_INV_1 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y78__R3_BUF_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y79__R0_BUF_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R0_INV_0 (.A(tie_lo_T0Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y79__R1_BUF_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R1_INV_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R2_INV_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y79__R2_INV_1 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y79__R3_BUF_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y7__R0_BUF_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R0_INV_0 (.A(tie_lo_T0Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y7__R1_BUF_0 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R1_INV_0 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R2_INV_0 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y7__R2_INV_1 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y7__R3_BUF_0 (.A(tie_lo_T0Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y80__R0_BUF_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R0_INV_0 (.A(tie_lo_T0Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y80__R1_BUF_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R1_INV_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R2_INV_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y80__R2_INV_1 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y80__R3_BUF_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y81__R0_BUF_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R0_INV_0 (.A(tie_lo_T0Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y81__R1_BUF_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R1_INV_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R2_INV_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y81__R2_INV_1 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y81__R3_BUF_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y82__R0_BUF_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R0_INV_0 (.A(tie_lo_T0Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y82__R1_BUF_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R1_INV_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R2_INV_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y82__R2_INV_1 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y82__R3_BUF_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y83__R0_BUF_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R0_INV_0 (.A(tie_lo_T0Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y83__R1_BUF_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R1_INV_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R2_INV_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y83__R2_INV_1 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y83__R3_BUF_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y84__R0_BUF_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R0_INV_0 (.A(tie_lo_T0Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y84__R1_BUF_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R1_INV_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R2_INV_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y84__R2_INV_1 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y84__R3_BUF_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y85__R0_BUF_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R0_INV_0 (.A(tie_lo_T0Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y85__R1_BUF_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R1_INV_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R2_INV_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y85__R2_INV_1 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y85__R3_BUF_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y86__R0_BUF_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R0_INV_0 (.A(tie_lo_T0Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y86__R1_BUF_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R1_INV_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R2_INV_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y86__R2_INV_1 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y86__R3_BUF_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y87__R0_BUF_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R0_INV_0 (.A(tie_lo_T0Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y87__R1_BUF_0 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R1_INV_0 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R2_INV_0 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y87__R2_INV_1 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y87__R3_BUF_0 (.A(tie_lo_T0Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y88__R0_BUF_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R0_INV_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y88__R1_BUF_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R1_INV_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R2_INV_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y88__R2_INV_1 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y88__R3_BUF_0 (.A(tie_lo_T0Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y89__R0_BUF_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R0_INV_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y89__R1_BUF_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R1_INV_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R2_INV_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y89__R2_INV_1 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y89__R3_BUF_0 (.A(tie_lo_T0Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y8__R0_BUF_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R0_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y8__R1_BUF_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R1_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R2_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y8__R2_INV_1 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y8__R3_BUF_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y9__R0_BUF_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R0_INV_0 (.A(tie_lo_T0Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y9__R1_BUF_0 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R1_INV_0 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T0Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R2_INV_0 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T0Y9__R2_INV_1 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T0Y9__R3_BUF_0 (.A(tie_lo_T0Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y0__R0_BUF_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R0_INV_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y0__R1_BUF_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R1_INV_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R2_INV_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y0__R2_INV_1 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y0__R3_BUF_0 (.A(tie_lo_T10Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y10__R0_BUF_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R0_INV_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y10__R1_BUF_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R1_INV_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R2_INV_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y10__R2_INV_1 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y10__R3_BUF_0 (.A(tie_lo_T10Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y11__R0_BUF_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R0_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y11__R1_BUF_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R1_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R2_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y11__R2_INV_1 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y11__R3_BUF_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y12__R0_BUF_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R0_INV_0 (.A(tie_lo_T10Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y12__R1_BUF_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R1_INV_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R2_INV_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y12__R2_INV_1 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y12__R3_BUF_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y13__R0_BUF_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R0_INV_0 (.A(tie_lo_T10Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y13__R1_BUF_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R1_INV_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R2_INV_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y13__R2_INV_1 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y13__R3_BUF_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y14__R0_BUF_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R0_INV_0 (.A(tie_lo_T10Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y14__R1_BUF_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R1_INV_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R2_INV_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y14__R2_INV_1 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y14__R3_BUF_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y15__R0_BUF_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R0_INV_0 (.A(tie_lo_T10Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y15__R1_BUF_0 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R1_INV_0 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R2_INV_0 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y15__R2_INV_1 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y15__R3_BUF_0 (.A(tie_lo_T10Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y16__R0_BUF_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R0_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y16__R1_BUF_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R1_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R2_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y16__R2_INV_1 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y16__R3_BUF_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y17__R0_BUF_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R0_INV_0 (.A(tie_lo_T10Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y17__R1_BUF_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R1_INV_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R2_INV_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y17__R2_INV_1 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y17__R3_BUF_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y18__R0_BUF_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R0_INV_0 (.A(tie_lo_T10Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y18__R1_BUF_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R1_INV_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R2_INV_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y18__R2_INV_1 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y18__R3_BUF_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y19__R0_BUF_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R0_INV_0 (.A(tie_lo_T10Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y19__R1_BUF_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R1_INV_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R2_INV_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y19__R2_INV_1 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y19__R3_BUF_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y1__R0_BUF_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R0_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y1__R1_BUF_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R1_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R2_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y1__R2_INV_1 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y1__R3_BUF_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y20__R0_BUF_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R0_INV_0 (.A(tie_lo_T10Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y20__R1_BUF_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R1_INV_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R2_INV_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y20__R2_INV_1 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y20__R3_BUF_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y21__R0_BUF_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R0_INV_0 (.A(tie_lo_T10Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y21__R1_BUF_0 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R1_INV_0 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R2_INV_0 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y21__R2_INV_1 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y21__R3_BUF_0 (.A(tie_lo_T10Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y22__R0_BUF_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R0_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y22__R1_BUF_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R1_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R2_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y22__R2_INV_1 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y22__R3_BUF_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y23__R0_BUF_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R0_INV_0 (.A(tie_lo_T10Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y23__R1_BUF_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R1_INV_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R2_INV_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y23__R2_INV_1 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y23__R3_BUF_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y24__R0_BUF_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R0_INV_0 (.A(tie_lo_T10Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y24__R1_BUF_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R1_INV_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R2_INV_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y24__R2_INV_1 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y24__R3_BUF_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y25__R0_BUF_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R0_INV_0 (.A(tie_lo_T10Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y25__R1_BUF_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R1_INV_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R2_INV_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y25__R2_INV_1 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y25__R3_BUF_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y26__R0_BUF_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R0_INV_0 (.A(tie_lo_T10Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y26__R1_BUF_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R1_INV_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R2_INV_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y26__R2_INV_1 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y26__R3_BUF_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y27__R0_BUF_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R0_INV_0 (.A(tie_lo_T10Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y27__R1_BUF_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R1_INV_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R2_INV_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y27__R2_INV_1 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y27__R3_BUF_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y28__R0_BUF_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R0_INV_0 (.A(tie_lo_T10Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y28__R1_BUF_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R1_INV_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R2_INV_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y28__R2_INV_1 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y28__R3_BUF_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y29__R0_BUF_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R0_INV_0 (.A(tie_lo_T10Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y29__R1_BUF_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R1_INV_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R2_INV_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y29__R2_INV_1 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y29__R3_BUF_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y2__R0_BUF_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R0_INV_0 (.A(tie_lo_T10Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y2__R1_BUF_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R1_INV_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R2_INV_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y2__R2_INV_1 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y2__R3_BUF_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y30__R0_BUF_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R0_INV_0 (.A(tie_lo_T10Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y30__R1_BUF_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R1_INV_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R2_INV_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y30__R2_INV_1 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y30__R3_BUF_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y31__R0_BUF_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R0_INV_0 (.A(tie_lo_T10Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y31__R1_BUF_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R1_INV_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R2_INV_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y31__R2_INV_1 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y31__R3_BUF_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y32__R0_BUF_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R0_INV_0 (.A(tie_lo_T10Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y32__R1_BUF_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R1_INV_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R2_INV_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y32__R2_INV_1 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y32__R3_BUF_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y33__R0_BUF_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R0_INV_0 (.A(tie_lo_T10Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y33__R1_BUF_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R1_INV_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R2_INV_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y33__R2_INV_1 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y33__R3_BUF_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y34__R0_BUF_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R0_INV_0 (.A(tie_lo_T10Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y34__R1_BUF_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R1_INV_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R2_INV_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y34__R2_INV_1 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y34__R3_BUF_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y35__R0_BUF_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R0_INV_0 (.A(tie_lo_T10Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y35__R1_BUF_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R1_INV_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R2_INV_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y35__R2_INV_1 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y35__R3_BUF_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y36__R0_BUF_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R0_INV_0 (.A(tie_lo_T10Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y36__R1_BUF_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R1_INV_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R2_INV_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y36__R2_INV_1 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y36__R3_BUF_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y37__R0_BUF_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R0_INV_0 (.A(tie_lo_T10Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y37__R1_BUF_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R1_INV_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R2_INV_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y37__R2_INV_1 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y37__R3_BUF_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y38__R0_BUF_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R0_INV_0 (.A(tie_lo_T10Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y38__R1_BUF_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R1_INV_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R2_INV_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y38__R2_INV_1 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y38__R3_BUF_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y39__R0_BUF_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R0_INV_0 (.A(tie_lo_T10Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y39__R1_BUF_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R1_INV_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R2_INV_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y39__R2_INV_1 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y39__R3_BUF_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y3__R0_BUF_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R0_INV_0 (.A(tie_lo_T10Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y3__R1_BUF_0 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R1_INV_0 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R2_INV_0 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y3__R2_INV_1 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y3__R3_BUF_0 (.A(tie_lo_T10Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y40__R0_BUF_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R0_INV_0 (.A(tie_lo_T10Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y40__R1_BUF_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R1_INV_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R2_INV_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y40__R2_INV_1 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y40__R3_BUF_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y41__R0_BUF_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R0_INV_0 (.A(tie_lo_T10Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y41__R1_BUF_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R1_INV_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R2_INV_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y41__R2_INV_1 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y41__R3_BUF_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y42__R0_BUF_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R0_INV_0 (.A(tie_lo_T10Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y42__R1_BUF_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R1_INV_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R2_INV_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y42__R2_INV_1 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y42__R3_BUF_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y43__R0_BUF_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R0_INV_0 (.A(tie_lo_T10Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y43__R1_BUF_0 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R1_INV_0 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R2_INV_0 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y43__R2_INV_1 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y43__R3_BUF_0 (.A(tie_lo_T10Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y44__R0_BUF_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R0_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y44__R1_BUF_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R1_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R2_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y44__R2_INV_1 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y44__R3_BUF_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y45__R0_BUF_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R0_INV_0 (.A(tie_lo_T10Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y45__R1_BUF_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R1_INV_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R2_INV_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y45__R2_INV_1 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y45__R3_BUF_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y46__R0_BUF_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R0_INV_0 (.A(tie_lo_T10Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y46__R1_BUF_0 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R1_INV_0 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R2_INV_0 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y46__R2_INV_1 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y46__R3_BUF_0 (.A(tie_lo_T10Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y47__R0_BUF_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R0_INV_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y47__R1_BUF_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R1_INV_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R2_INV_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y47__R2_INV_1 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y47__R3_BUF_0 (.A(tie_lo_T10Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y48__R0_BUF_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R0_INV_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y48__R1_BUF_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R1_INV_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R2_INV_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y48__R2_INV_1 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y48__R3_BUF_0 (.A(tie_lo_T10Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y49__R0_BUF_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R0_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y49__R1_BUF_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R1_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R2_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y49__R2_INV_1 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y49__R3_BUF_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y4__R0_BUF_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R0_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y4__R1_BUF_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R1_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R2_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y4__R2_INV_1 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y4__R3_BUF_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y50__R0_BUF_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R0_INV_0 (.A(tie_lo_T10Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y50__R1_BUF_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R1_INV_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R2_INV_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y50__R2_INV_1 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y50__R3_BUF_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y51__R0_BUF_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R0_INV_0 (.A(tie_lo_T10Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y51__R1_BUF_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R1_INV_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R2_INV_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y51__R2_INV_1 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y51__R3_BUF_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y52__R0_BUF_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R0_INV_0 (.A(tie_lo_T10Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y52__R1_BUF_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R1_INV_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R2_INV_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y52__R2_INV_1 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y52__R3_BUF_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y53__R0_BUF_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R0_INV_0 (.A(tie_lo_T10Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y53__R1_BUF_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R1_INV_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R2_INV_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y53__R2_INV_1 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y53__R3_BUF_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y54__R0_BUF_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R0_INV_0 (.A(tie_lo_T10Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y54__R1_BUF_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R1_INV_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R2_INV_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y54__R2_INV_1 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y54__R3_BUF_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y55__R0_BUF_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R0_INV_0 (.A(tie_lo_T10Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y55__R1_BUF_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R1_INV_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R2_INV_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y55__R2_INV_1 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y55__R3_BUF_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y56__R0_BUF_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R0_INV_0 (.A(tie_lo_T10Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y56__R1_BUF_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R1_INV_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R2_INV_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y56__R2_INV_1 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y56__R3_BUF_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y57__R0_BUF_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R0_INV_0 (.A(tie_lo_T10Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y57__R1_BUF_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R1_INV_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R2_INV_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y57__R2_INV_1 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y57__R3_BUF_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y58__R0_BUF_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R0_INV_0 (.A(tie_lo_T10Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y58__R1_BUF_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R1_INV_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R2_INV_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y58__R2_INV_1 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y58__R3_BUF_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y59__R0_BUF_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R0_INV_0 (.A(tie_lo_T10Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y59__R1_BUF_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R1_INV_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R2_INV_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y59__R2_INV_1 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y59__R3_BUF_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y5__R0_BUF_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R0_INV_0 (.A(tie_lo_T10Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y5__R1_BUF_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R1_INV_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R2_INV_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y5__R2_INV_1 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y5__R3_BUF_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y60__R0_BUF_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R0_INV_0 (.A(tie_lo_T10Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y60__R1_BUF_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R1_INV_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R2_INV_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y60__R2_INV_1 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y60__R3_BUF_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y61__R0_BUF_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R0_INV_0 (.A(tie_lo_T10Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y61__R1_BUF_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R1_INV_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R2_INV_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y61__R2_INV_1 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y61__R3_BUF_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y62__R0_BUF_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R0_INV_0 (.A(tie_lo_T10Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y62__R1_BUF_0 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R1_INV_0 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R2_INV_0 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y62__R2_INV_1 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y62__R3_BUF_0 (.A(tie_lo_T10Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y63__R0_BUF_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R0_INV_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y63__R1_BUF_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R1_INV_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R2_INV_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y63__R2_INV_1 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y63__R3_BUF_0 (.A(tie_lo_T10Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y64__R0_BUF_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R0_INV_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y64__R1_BUF_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R1_INV_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R2_INV_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y64__R2_INV_1 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y64__R3_BUF_0 (.A(tie_lo_T10Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y65__R0_BUF_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R0_INV_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y65__R1_BUF_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R1_INV_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R2_INV_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y65__R2_INV_1 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y65__R3_BUF_0 (.A(tie_lo_T10Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y66__R0_BUF_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R0_INV_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y66__R1_BUF_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R1_INV_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R2_INV_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y66__R2_INV_1 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y66__R3_BUF_0 (.A(tie_lo_T10Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y67__R0_BUF_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R0_INV_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y67__R1_BUF_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R1_INV_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R2_INV_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y67__R2_INV_1 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y67__R3_BUF_0 (.A(tie_lo_T10Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y68__R0_BUF_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R0_INV_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y68__R1_BUF_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R1_INV_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R2_INV_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y68__R2_INV_1 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y68__R3_BUF_0 (.A(tie_lo_T10Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y69__R0_BUF_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R0_INV_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y69__R1_BUF_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R1_INV_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R2_INV_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y69__R2_INV_1 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y69__R3_BUF_0 (.A(tie_lo_T10Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y6__R0_BUF_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R0_INV_0 (.A(tie_lo_T10Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y6__R1_BUF_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R1_INV_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R2_INV_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y6__R2_INV_1 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y6__R3_BUF_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y70__R0_BUF_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R0_INV_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y70__R1_BUF_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R1_INV_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R2_INV_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y70__R2_INV_1 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y70__R3_BUF_0 (.A(tie_lo_T10Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y71__R0_BUF_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R0_INV_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y71__R1_BUF_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R1_INV_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R2_INV_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y71__R2_INV_1 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y71__R3_BUF_0 (.A(tie_lo_T10Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y72__R0_BUF_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R0_INV_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y72__R1_BUF_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R1_INV_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R2_INV_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y72__R2_INV_1 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y72__R3_BUF_0 (.A(tie_lo_T10Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y73__R0_BUF_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R0_INV_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y73__R1_BUF_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R1_INV_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R2_INV_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y73__R2_INV_1 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y73__R3_BUF_0 (.A(tie_lo_T10Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y74__R0_BUF_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R0_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y74__R1_BUF_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R1_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R2_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y74__R2_INV_1 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y74__R3_BUF_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y75__R0_BUF_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R0_INV_0 (.A(tie_lo_T10Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y75__R1_BUF_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R1_INV_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R2_INV_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y75__R2_INV_1 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y75__R3_BUF_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y76__R0_BUF_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R0_INV_0 (.A(tie_lo_T10Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y76__R1_BUF_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R1_INV_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R2_INV_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y76__R2_INV_1 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y76__R3_BUF_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y77__R0_BUF_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R0_INV_0 (.A(tie_lo_T10Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y77__R1_BUF_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R1_INV_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R2_INV_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y77__R2_INV_1 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y77__R3_BUF_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y78__R0_BUF_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R0_INV_0 (.A(tie_lo_T10Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y78__R1_BUF_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R1_INV_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R2_INV_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y78__R2_INV_1 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y78__R3_BUF_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y79__R0_BUF_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R0_INV_0 (.A(tie_lo_T10Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y79__R1_BUF_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R1_INV_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R2_INV_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y79__R2_INV_1 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y79__R3_BUF_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y7__R0_BUF_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R0_INV_0 (.A(tie_lo_T10Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y7__R1_BUF_0 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R1_INV_0 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R2_INV_0 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y7__R2_INV_1 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y7__R3_BUF_0 (.A(tie_lo_T10Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y80__R0_BUF_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R0_INV_0 (.A(tie_lo_T10Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y80__R1_BUF_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R1_INV_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R2_INV_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y80__R2_INV_1 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y80__R3_BUF_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y81__R0_BUF_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R0_INV_0 (.A(tie_lo_T10Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y81__R1_BUF_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R1_INV_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R2_INV_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y81__R2_INV_1 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y81__R3_BUF_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y82__R0_BUF_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R0_INV_0 (.A(tie_lo_T10Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y82__R1_BUF_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R1_INV_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R2_INV_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y82__R2_INV_1 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y82__R3_BUF_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y83__R0_BUF_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R0_INV_0 (.A(tie_lo_T10Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y83__R1_BUF_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R1_INV_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R2_INV_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y83__R2_INV_1 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y83__R3_BUF_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y84__R0_BUF_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R0_INV_0 (.A(tie_lo_T10Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y84__R1_BUF_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R1_INV_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R2_INV_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y84__R2_INV_1 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y84__R3_BUF_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y85__R0_BUF_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R0_INV_0 (.A(tie_lo_T10Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y85__R1_BUF_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R1_INV_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R2_INV_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y85__R2_INV_1 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y85__R3_BUF_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y86__R0_BUF_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R0_INV_0 (.A(tie_lo_T10Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y86__R1_BUF_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R1_INV_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R2_INV_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y86__R2_INV_1 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y86__R3_BUF_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y87__R0_BUF_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R0_INV_0 (.A(tie_lo_T10Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y87__R1_BUF_0 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R1_INV_0 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R2_INV_0 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y87__R2_INV_1 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y87__R3_BUF_0 (.A(tie_lo_T10Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y88__R0_BUF_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R0_INV_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y88__R1_BUF_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R1_INV_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R2_INV_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y88__R2_INV_1 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y88__R3_BUF_0 (.A(tie_lo_T10Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y89__R0_BUF_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R0_INV_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y89__R1_BUF_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R1_INV_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R2_INV_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y89__R2_INV_1 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y89__R3_BUF_0 (.A(tie_lo_T10Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y8__R0_BUF_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R0_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y8__R1_BUF_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R1_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R2_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y8__R2_INV_1 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y8__R3_BUF_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y9__R0_BUF_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R0_INV_0 (.A(tie_lo_T10Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y9__R1_BUF_0 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R1_INV_0 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T10Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R2_INV_0 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T10Y9__R2_INV_1 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T10Y9__R3_BUF_0 (.A(tie_lo_T10Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y0__R0_BUF_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R0_INV_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y0__R1_BUF_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R1_INV_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R2_INV_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y0__R2_INV_1 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y0__R3_BUF_0 (.A(tie_lo_T11Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y10__R0_BUF_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R0_INV_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y10__R1_BUF_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R1_INV_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R2_INV_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y10__R2_INV_1 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y10__R3_BUF_0 (.A(tie_lo_T11Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y11__R0_BUF_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R0_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y11__R1_BUF_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R1_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R2_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y11__R2_INV_1 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y11__R3_BUF_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y12__R0_BUF_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R0_INV_0 (.A(tie_lo_T11Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y12__R1_BUF_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R1_INV_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R2_INV_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y12__R2_INV_1 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y12__R3_BUF_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y13__R0_BUF_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R0_INV_0 (.A(tie_lo_T11Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y13__R1_BUF_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R1_INV_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R2_INV_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y13__R2_INV_1 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y13__R3_BUF_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y14__R0_BUF_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R0_INV_0 (.A(tie_lo_T11Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y14__R1_BUF_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R1_INV_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R2_INV_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y14__R2_INV_1 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y14__R3_BUF_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y15__R0_BUF_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R0_INV_0 (.A(tie_lo_T11Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y15__R1_BUF_0 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R1_INV_0 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R2_INV_0 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y15__R2_INV_1 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y15__R3_BUF_0 (.A(tie_lo_T11Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y16__R0_BUF_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R0_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y16__R1_BUF_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R1_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R2_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y16__R2_INV_1 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y16__R3_BUF_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y17__R0_BUF_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R0_INV_0 (.A(tie_lo_T11Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y17__R1_BUF_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R1_INV_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R2_INV_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y17__R2_INV_1 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y17__R3_BUF_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y18__R0_BUF_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R0_INV_0 (.A(tie_lo_T11Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y18__R1_BUF_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R1_INV_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R2_INV_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y18__R2_INV_1 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y18__R3_BUF_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y19__R0_BUF_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R0_INV_0 (.A(tie_lo_T11Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y19__R1_BUF_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R1_INV_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R2_INV_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y19__R2_INV_1 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y19__R3_BUF_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y1__R0_BUF_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R0_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y1__R1_BUF_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R1_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R2_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y1__R2_INV_1 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y1__R3_BUF_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y20__R0_BUF_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R0_INV_0 (.A(tie_lo_T11Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y20__R1_BUF_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R1_INV_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R2_INV_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y20__R2_INV_1 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y20__R3_BUF_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y21__R0_BUF_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R0_INV_0 (.A(tie_lo_T11Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y21__R1_BUF_0 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R1_INV_0 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R2_INV_0 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y21__R2_INV_1 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y21__R3_BUF_0 (.A(tie_lo_T11Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y22__R0_BUF_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R0_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y22__R1_BUF_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R1_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R2_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y22__R2_INV_1 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y22__R3_BUF_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y23__R0_BUF_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R0_INV_0 (.A(tie_lo_T11Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y23__R1_BUF_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R1_INV_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R2_INV_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y23__R2_INV_1 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y23__R3_BUF_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y24__R0_BUF_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R0_INV_0 (.A(tie_lo_T11Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y24__R1_BUF_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R1_INV_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R2_INV_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y24__R2_INV_1 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y24__R3_BUF_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y25__R0_BUF_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R0_INV_0 (.A(tie_lo_T11Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y25__R1_BUF_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R1_INV_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R2_INV_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y25__R2_INV_1 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y25__R3_BUF_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y26__R0_BUF_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R0_INV_0 (.A(tie_lo_T11Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y26__R1_BUF_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R1_INV_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R2_INV_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y26__R2_INV_1 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y26__R3_BUF_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y27__R0_BUF_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R0_INV_0 (.A(tie_lo_T11Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y27__R1_BUF_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R1_INV_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R2_INV_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y27__R2_INV_1 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y27__R3_BUF_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y28__R0_BUF_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R0_INV_0 (.A(tie_lo_T11Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y28__R1_BUF_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R1_INV_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R2_INV_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y28__R2_INV_1 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y28__R3_BUF_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y29__R0_BUF_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R0_INV_0 (.A(tie_lo_T11Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y29__R1_BUF_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R1_INV_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R2_INV_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y29__R2_INV_1 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y29__R3_BUF_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y2__R0_BUF_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R0_INV_0 (.A(tie_lo_T11Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y2__R1_BUF_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R1_INV_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R2_INV_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y2__R2_INV_1 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y2__R3_BUF_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y30__R0_BUF_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R0_INV_0 (.A(tie_lo_T11Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y30__R1_BUF_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R1_INV_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R2_INV_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y30__R2_INV_1 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y30__R3_BUF_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y31__R0_BUF_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R0_INV_0 (.A(tie_lo_T11Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y31__R1_BUF_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R1_INV_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R2_INV_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y31__R2_INV_1 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y31__R3_BUF_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y32__R0_BUF_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R0_INV_0 (.A(tie_lo_T11Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y32__R1_BUF_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R1_INV_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R2_INV_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y32__R2_INV_1 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y32__R3_BUF_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y33__R0_BUF_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R0_INV_0 (.A(tie_lo_T11Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y33__R1_BUF_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R1_INV_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R2_INV_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y33__R2_INV_1 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y33__R3_BUF_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y34__R0_BUF_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R0_INV_0 (.A(tie_lo_T11Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y34__R1_BUF_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R1_INV_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R2_INV_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y34__R2_INV_1 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y34__R3_BUF_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y35__R0_BUF_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R0_INV_0 (.A(tie_lo_T11Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y35__R1_BUF_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R1_INV_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R2_INV_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y35__R2_INV_1 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y35__R3_BUF_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y36__R0_BUF_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R0_INV_0 (.A(tie_lo_T11Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y36__R1_BUF_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R1_INV_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R2_INV_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y36__R2_INV_1 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y36__R3_BUF_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y37__R0_BUF_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R0_INV_0 (.A(tie_lo_T11Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y37__R1_BUF_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R1_INV_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R2_INV_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y37__R2_INV_1 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y37__R3_BUF_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y38__R0_BUF_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R0_INV_0 (.A(tie_lo_T11Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y38__R1_BUF_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R1_INV_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R2_INV_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y38__R2_INV_1 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y38__R3_BUF_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y39__R0_BUF_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R0_INV_0 (.A(tie_lo_T11Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y39__R1_BUF_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R1_INV_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R2_INV_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y39__R2_INV_1 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y39__R3_BUF_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y3__R0_BUF_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R0_INV_0 (.A(tie_lo_T11Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y3__R1_BUF_0 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R1_INV_0 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R2_INV_0 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y3__R2_INV_1 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y3__R3_BUF_0 (.A(tie_lo_T11Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y40__R0_BUF_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R0_INV_0 (.A(tie_lo_T11Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y40__R1_BUF_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R1_INV_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R2_INV_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y40__R2_INV_1 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y40__R3_BUF_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y41__R0_BUF_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R0_INV_0 (.A(tie_lo_T11Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y41__R1_BUF_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R1_INV_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R2_INV_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y41__R2_INV_1 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y41__R3_BUF_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y42__R0_BUF_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R0_INV_0 (.A(tie_lo_T11Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y42__R1_BUF_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R1_INV_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R2_INV_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y42__R2_INV_1 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y42__R3_BUF_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y43__R0_BUF_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R0_INV_0 (.A(tie_lo_T11Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y43__R1_BUF_0 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R1_INV_0 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R2_INV_0 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y43__R2_INV_1 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y43__R3_BUF_0 (.A(tie_lo_T11Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y44__R0_BUF_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R0_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y44__R1_BUF_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R1_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R2_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y44__R2_INV_1 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y44__R3_BUF_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y45__R0_BUF_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R0_INV_0 (.A(tie_lo_T11Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y45__R1_BUF_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R1_INV_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R2_INV_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y45__R2_INV_1 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y45__R3_BUF_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y46__R0_BUF_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R0_INV_0 (.A(tie_lo_T11Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y46__R1_BUF_0 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R1_INV_0 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R2_INV_0 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y46__R2_INV_1 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y46__R3_BUF_0 (.A(tie_lo_T11Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y47__R0_BUF_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R0_INV_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y47__R1_BUF_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R1_INV_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R2_INV_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y47__R2_INV_1 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y47__R3_BUF_0 (.A(tie_lo_T11Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y48__R0_BUF_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R0_INV_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y48__R1_BUF_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R1_INV_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R2_INV_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y48__R2_INV_1 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y48__R3_BUF_0 (.A(tie_lo_T11Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y49__R0_BUF_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R0_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y49__R1_BUF_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R1_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R2_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y49__R2_INV_1 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y49__R3_BUF_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y4__R0_BUF_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R0_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y4__R1_BUF_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R1_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R2_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y4__R2_INV_1 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y4__R3_BUF_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y50__R0_BUF_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R0_INV_0 (.A(tie_lo_T11Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y50__R1_BUF_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R1_INV_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R2_INV_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y50__R2_INV_1 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y50__R3_BUF_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y51__R0_BUF_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R0_INV_0 (.A(tie_lo_T11Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y51__R1_BUF_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R1_INV_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R2_INV_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y51__R2_INV_1 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y51__R3_BUF_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y52__R0_BUF_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R0_INV_0 (.A(tie_lo_T11Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y52__R1_BUF_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R1_INV_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R2_INV_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y52__R2_INV_1 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y52__R3_BUF_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y53__R0_BUF_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R0_INV_0 (.A(tie_lo_T11Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y53__R1_BUF_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R1_INV_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R2_INV_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y53__R2_INV_1 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y53__R3_BUF_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y54__R0_BUF_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R0_INV_0 (.A(tie_lo_T11Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y54__R1_BUF_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R1_INV_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R2_INV_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y54__R2_INV_1 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y54__R3_BUF_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y55__R0_BUF_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R0_INV_0 (.A(tie_lo_T11Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y55__R1_BUF_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R1_INV_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R2_INV_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y55__R2_INV_1 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y55__R3_BUF_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y56__R0_BUF_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R0_INV_0 (.A(tie_lo_T11Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y56__R1_BUF_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R1_INV_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R2_INV_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y56__R2_INV_1 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y56__R3_BUF_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y57__R0_BUF_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R0_INV_0 (.A(tie_lo_T11Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y57__R1_BUF_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R1_INV_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R2_INV_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y57__R2_INV_1 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y57__R3_BUF_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y58__R0_BUF_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R0_INV_0 (.A(tie_lo_T11Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y58__R1_BUF_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R1_INV_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R2_INV_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y58__R2_INV_1 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y58__R3_BUF_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y59__R0_BUF_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R0_INV_0 (.A(tie_lo_T11Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y59__R1_BUF_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R1_INV_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R2_INV_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y59__R2_INV_1 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y59__R3_BUF_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y5__R0_BUF_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R0_INV_0 (.A(tie_lo_T11Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y5__R1_BUF_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R1_INV_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R2_INV_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y5__R2_INV_1 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y5__R3_BUF_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y60__R0_BUF_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R0_INV_0 (.A(tie_lo_T11Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y60__R1_BUF_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R1_INV_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R2_INV_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y60__R2_INV_1 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y60__R3_BUF_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y61__R0_BUF_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R0_INV_0 (.A(tie_lo_T11Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y61__R1_BUF_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R1_INV_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R2_INV_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y61__R2_INV_1 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y61__R3_BUF_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y62__R0_BUF_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R0_INV_0 (.A(tie_lo_T11Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y62__R1_BUF_0 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R1_INV_0 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R2_INV_0 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y62__R2_INV_1 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y62__R3_BUF_0 (.A(tie_lo_T11Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y63__R0_BUF_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R0_INV_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y63__R1_BUF_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R1_INV_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R2_INV_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y63__R2_INV_1 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y63__R3_BUF_0 (.A(tie_lo_T11Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y64__R0_BUF_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R0_INV_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y64__R1_BUF_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R1_INV_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R2_INV_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y64__R2_INV_1 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y64__R3_BUF_0 (.A(tie_lo_T11Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y65__R0_BUF_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R0_INV_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y65__R1_BUF_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R1_INV_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R2_INV_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y65__R2_INV_1 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y65__R3_BUF_0 (.A(tie_lo_T11Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y66__R0_BUF_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R0_INV_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y66__R1_BUF_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R1_INV_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R2_INV_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y66__R2_INV_1 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y66__R3_BUF_0 (.A(tie_lo_T11Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y67__R0_BUF_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R0_INV_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y67__R1_BUF_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R1_INV_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R2_INV_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y67__R2_INV_1 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y67__R3_BUF_0 (.A(tie_lo_T11Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y68__R0_BUF_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R0_INV_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y68__R1_BUF_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R1_INV_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R2_INV_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y68__R2_INV_1 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y68__R3_BUF_0 (.A(tie_lo_T11Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y69__R0_BUF_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R0_INV_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y69__R1_BUF_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R1_INV_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R2_INV_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y69__R2_INV_1 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y69__R3_BUF_0 (.A(tie_lo_T11Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y6__R0_BUF_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R0_INV_0 (.A(tie_lo_T11Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y6__R1_BUF_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R1_INV_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R2_INV_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y6__R2_INV_1 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y6__R3_BUF_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y70__R0_BUF_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R0_INV_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y70__R1_BUF_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R1_INV_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R2_INV_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y70__R2_INV_1 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y70__R3_BUF_0 (.A(tie_lo_T11Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y71__R0_BUF_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R0_INV_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y71__R1_BUF_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R1_INV_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R2_INV_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y71__R2_INV_1 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y71__R3_BUF_0 (.A(tie_lo_T11Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y72__R0_BUF_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R0_INV_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y72__R1_BUF_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R1_INV_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R2_INV_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y72__R2_INV_1 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y72__R3_BUF_0 (.A(tie_lo_T11Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y73__R0_BUF_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R0_INV_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y73__R1_BUF_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R1_INV_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R2_INV_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y73__R2_INV_1 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y73__R3_BUF_0 (.A(tie_lo_T11Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y74__R0_BUF_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R0_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y74__R1_BUF_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R1_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R2_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y74__R2_INV_1 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y74__R3_BUF_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y75__R0_BUF_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R0_INV_0 (.A(tie_lo_T11Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y75__R1_BUF_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R1_INV_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R2_INV_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y75__R2_INV_1 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y75__R3_BUF_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y76__R0_BUF_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R0_INV_0 (.A(tie_lo_T11Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y76__R1_BUF_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R1_INV_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R2_INV_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y76__R2_INV_1 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y76__R3_BUF_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y77__R0_BUF_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R0_INV_0 (.A(tie_lo_T11Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y77__R1_BUF_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R1_INV_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R2_INV_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y77__R2_INV_1 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y77__R3_BUF_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y78__R0_BUF_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R0_INV_0 (.A(tie_lo_T11Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y78__R1_BUF_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R1_INV_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R2_INV_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y78__R2_INV_1 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y78__R3_BUF_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y79__R0_BUF_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R0_INV_0 (.A(tie_lo_T11Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y79__R1_BUF_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R1_INV_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R2_INV_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y79__R2_INV_1 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y79__R3_BUF_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y7__R0_BUF_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R0_INV_0 (.A(tie_lo_T11Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y7__R1_BUF_0 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R1_INV_0 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R2_INV_0 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y7__R2_INV_1 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y7__R3_BUF_0 (.A(tie_lo_T11Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y80__R0_BUF_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R0_INV_0 (.A(tie_lo_T11Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y80__R1_BUF_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R1_INV_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R2_INV_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y80__R2_INV_1 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y80__R3_BUF_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y81__R0_BUF_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R0_INV_0 (.A(tie_lo_T11Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y81__R1_BUF_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R1_INV_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R2_INV_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y81__R2_INV_1 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y81__R3_BUF_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y82__R0_BUF_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R0_INV_0 (.A(tie_lo_T11Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y82__R1_BUF_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R1_INV_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R2_INV_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y82__R2_INV_1 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y82__R3_BUF_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y83__R0_BUF_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R0_INV_0 (.A(tie_lo_T11Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y83__R1_BUF_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R1_INV_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R2_INV_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y83__R2_INV_1 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y83__R3_BUF_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y84__R0_BUF_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R0_INV_0 (.A(tie_lo_T11Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y84__R1_BUF_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R1_INV_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R2_INV_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y84__R2_INV_1 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y84__R3_BUF_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y85__R0_BUF_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R0_INV_0 (.A(tie_lo_T11Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y85__R1_BUF_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R1_INV_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R2_INV_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y85__R2_INV_1 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y85__R3_BUF_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y86__R0_BUF_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R0_INV_0 (.A(tie_lo_T11Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y86__R1_BUF_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R1_INV_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R2_INV_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y86__R2_INV_1 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y86__R3_BUF_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y87__R0_BUF_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R0_INV_0 (.A(tie_lo_T11Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y87__R1_BUF_0 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R1_INV_0 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R2_INV_0 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y87__R2_INV_1 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y87__R3_BUF_0 (.A(tie_lo_T11Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y88__R0_BUF_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R0_INV_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y88__R1_BUF_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R1_INV_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R2_INV_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y88__R2_INV_1 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y88__R3_BUF_0 (.A(tie_lo_T11Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y89__R0_BUF_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R0_INV_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y89__R1_BUF_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R1_INV_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R2_INV_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y89__R2_INV_1 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y89__R3_BUF_0 (.A(tie_lo_T11Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y8__R0_BUF_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R0_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y8__R1_BUF_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R1_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R2_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y8__R2_INV_1 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y8__R3_BUF_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y9__R0_BUF_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R0_INV_0 (.A(tie_lo_T11Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y9__R1_BUF_0 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R1_INV_0 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T11Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R2_INV_0 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T11Y9__R2_INV_1 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T11Y9__R3_BUF_0 (.A(tie_lo_T11Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y0__R0_BUF_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R0_INV_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y0__R1_BUF_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R1_INV_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R2_INV_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y0__R2_INV_1 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y0__R3_BUF_0 (.A(tie_lo_T12Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y10__R0_BUF_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R0_INV_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y10__R1_BUF_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R1_INV_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R2_INV_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y10__R2_INV_1 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y10__R3_BUF_0 (.A(tie_lo_T12Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y11__R0_BUF_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R0_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y11__R1_BUF_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R1_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R2_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y11__R2_INV_1 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y11__R3_BUF_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y12__R0_BUF_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R0_INV_0 (.A(tie_lo_T12Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y12__R1_BUF_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R1_INV_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R2_INV_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y12__R2_INV_1 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y12__R3_BUF_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y13__R0_BUF_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R0_INV_0 (.A(tie_lo_T12Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y13__R1_BUF_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R1_INV_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R2_INV_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y13__R2_INV_1 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y13__R3_BUF_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y14__R0_BUF_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R0_INV_0 (.A(tie_lo_T12Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y14__R1_BUF_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R1_INV_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R2_INV_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y14__R2_INV_1 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y14__R3_BUF_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y15__R0_BUF_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R0_INV_0 (.A(tie_lo_T12Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y15__R1_BUF_0 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R1_INV_0 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R2_INV_0 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y15__R2_INV_1 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y15__R3_BUF_0 (.A(tie_lo_T12Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y16__R0_BUF_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R0_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y16__R1_BUF_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R1_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R2_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y16__R2_INV_1 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y16__R3_BUF_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y17__R0_BUF_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R0_INV_0 (.A(tie_lo_T12Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y17__R1_BUF_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R1_INV_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R2_INV_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y17__R2_INV_1 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y17__R3_BUF_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y18__R0_BUF_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R0_INV_0 (.A(tie_lo_T12Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y18__R1_BUF_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R1_INV_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R2_INV_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y18__R2_INV_1 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y18__R3_BUF_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y19__R0_BUF_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R0_INV_0 (.A(tie_lo_T12Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y19__R1_BUF_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R1_INV_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R2_INV_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y19__R2_INV_1 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y19__R3_BUF_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y1__R0_BUF_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R0_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y1__R1_BUF_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R1_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R2_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y1__R2_INV_1 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y1__R3_BUF_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y20__R0_BUF_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R0_INV_0 (.A(tie_lo_T12Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y20__R1_BUF_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R1_INV_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R2_INV_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y20__R2_INV_1 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y20__R3_BUF_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y21__R0_BUF_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R0_INV_0 (.A(tie_lo_T12Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y21__R1_BUF_0 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R1_INV_0 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R2_INV_0 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y21__R2_INV_1 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y21__R3_BUF_0 (.A(tie_lo_T12Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y22__R0_BUF_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R0_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y22__R1_BUF_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R1_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R2_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y22__R2_INV_1 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y22__R3_BUF_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y23__R0_BUF_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R0_INV_0 (.A(tie_lo_T12Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y23__R1_BUF_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R1_INV_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R2_INV_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y23__R2_INV_1 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y23__R3_BUF_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y24__R0_BUF_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R0_INV_0 (.A(tie_lo_T12Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y24__R1_BUF_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R1_INV_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R2_INV_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y24__R2_INV_1 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y24__R3_BUF_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y25__R0_BUF_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R0_INV_0 (.A(tie_lo_T12Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y25__R1_BUF_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R1_INV_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R2_INV_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y25__R2_INV_1 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y25__R3_BUF_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y26__R0_BUF_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R0_INV_0 (.A(tie_lo_T12Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y26__R1_BUF_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R1_INV_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R2_INV_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y26__R2_INV_1 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y26__R3_BUF_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y27__R0_BUF_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R0_INV_0 (.A(tie_lo_T12Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y27__R1_BUF_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R1_INV_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R2_INV_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y27__R2_INV_1 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y27__R3_BUF_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y28__R0_BUF_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R0_INV_0 (.A(tie_lo_T12Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y28__R1_BUF_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R1_INV_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R2_INV_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y28__R2_INV_1 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y28__R3_BUF_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y29__R0_BUF_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R0_INV_0 (.A(tie_lo_T12Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y29__R1_BUF_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R1_INV_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R2_INV_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y29__R2_INV_1 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y29__R3_BUF_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y2__R0_BUF_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R0_INV_0 (.A(tie_lo_T12Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y2__R1_BUF_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R1_INV_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R2_INV_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y2__R2_INV_1 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y2__R3_BUF_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y30__R0_BUF_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R0_INV_0 (.A(tie_lo_T12Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y30__R1_BUF_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R1_INV_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R2_INV_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y30__R2_INV_1 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y30__R3_BUF_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y31__R0_BUF_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R0_INV_0 (.A(tie_lo_T12Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y31__R1_BUF_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R1_INV_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R2_INV_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y31__R2_INV_1 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y31__R3_BUF_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y32__R0_BUF_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R0_INV_0 (.A(tie_lo_T12Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y32__R1_BUF_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R1_INV_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R2_INV_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y32__R2_INV_1 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y32__R3_BUF_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y33__R0_BUF_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R0_INV_0 (.A(tie_lo_T12Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y33__R1_BUF_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R1_INV_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R2_INV_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y33__R2_INV_1 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y33__R3_BUF_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y34__R0_BUF_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R0_INV_0 (.A(tie_lo_T12Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y34__R1_BUF_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R1_INV_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R2_INV_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y34__R2_INV_1 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y34__R3_BUF_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y35__R0_BUF_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R0_INV_0 (.A(tie_lo_T12Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y35__R1_BUF_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R1_INV_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R2_INV_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y35__R2_INV_1 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y35__R3_BUF_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y36__R0_BUF_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R0_INV_0 (.A(tie_lo_T12Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y36__R1_BUF_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R1_INV_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R2_INV_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y36__R2_INV_1 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y36__R3_BUF_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y37__R0_BUF_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R0_INV_0 (.A(tie_lo_T12Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y37__R1_BUF_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R1_INV_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R2_INV_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y37__R2_INV_1 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y37__R3_BUF_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y38__R0_BUF_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R0_INV_0 (.A(tie_lo_T12Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y38__R1_BUF_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R1_INV_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R2_INV_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y38__R2_INV_1 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y38__R3_BUF_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y39__R0_BUF_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R0_INV_0 (.A(tie_lo_T12Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y39__R1_BUF_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R1_INV_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R2_INV_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y39__R2_INV_1 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y39__R3_BUF_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y3__R0_BUF_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R0_INV_0 (.A(tie_lo_T12Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y3__R1_BUF_0 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R1_INV_0 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R2_INV_0 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y3__R2_INV_1 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y3__R3_BUF_0 (.A(tie_lo_T12Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y40__R0_BUF_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R0_INV_0 (.A(tie_lo_T12Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y40__R1_BUF_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R1_INV_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R2_INV_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y40__R2_INV_1 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y40__R3_BUF_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y41__R0_BUF_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R0_INV_0 (.A(tie_lo_T12Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y41__R1_BUF_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R1_INV_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R2_INV_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y41__R2_INV_1 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y41__R3_BUF_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y42__R0_BUF_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R0_INV_0 (.A(tie_lo_T12Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y42__R1_BUF_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R1_INV_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R2_INV_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y42__R2_INV_1 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y42__R3_BUF_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y43__R0_BUF_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R0_INV_0 (.A(tie_lo_T12Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y43__R1_BUF_0 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R1_INV_0 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R2_INV_0 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y43__R2_INV_1 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y43__R3_BUF_0 (.A(tie_lo_T12Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y44__R0_BUF_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R0_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y44__R1_BUF_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R1_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R2_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y44__R2_INV_1 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y44__R3_BUF_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y45__R0_BUF_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R0_INV_0 (.A(tie_lo_T12Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y45__R1_BUF_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R1_INV_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R2_INV_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y45__R2_INV_1 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y45__R3_BUF_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y46__R0_BUF_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R0_INV_0 (.A(tie_lo_T12Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y46__R1_BUF_0 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R1_INV_0 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R2_INV_0 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y46__R2_INV_1 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y46__R3_BUF_0 (.A(tie_lo_T12Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y47__R0_BUF_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R0_INV_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y47__R1_BUF_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R1_INV_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R2_INV_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y47__R2_INV_1 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y47__R3_BUF_0 (.A(tie_lo_T12Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y48__R0_BUF_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R0_INV_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y48__R1_BUF_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R1_INV_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R2_INV_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y48__R2_INV_1 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y48__R3_BUF_0 (.A(tie_lo_T12Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y49__R0_BUF_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R0_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y49__R1_BUF_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R1_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R2_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y49__R2_INV_1 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y49__R3_BUF_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y4__R0_BUF_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R0_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y4__R1_BUF_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R1_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R2_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y4__R2_INV_1 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y4__R3_BUF_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y50__R0_BUF_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R0_INV_0 (.A(tie_lo_T12Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y50__R1_BUF_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R1_INV_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R2_INV_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y50__R2_INV_1 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y50__R3_BUF_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y51__R0_BUF_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R0_INV_0 (.A(tie_lo_T12Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y51__R1_BUF_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R1_INV_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R2_INV_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y51__R2_INV_1 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y51__R3_BUF_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y52__R0_BUF_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R0_INV_0 (.A(tie_lo_T12Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y52__R1_BUF_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R1_INV_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R2_INV_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y52__R2_INV_1 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y52__R3_BUF_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y53__R0_BUF_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R0_INV_0 (.A(tie_lo_T12Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y53__R1_BUF_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R1_INV_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R2_INV_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y53__R2_INV_1 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y53__R3_BUF_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y54__R0_BUF_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R0_INV_0 (.A(tie_lo_T12Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y54__R1_BUF_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R1_INV_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R2_INV_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y54__R2_INV_1 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y54__R3_BUF_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y55__R0_BUF_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R0_INV_0 (.A(tie_lo_T12Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y55__R1_BUF_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R1_INV_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R2_INV_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y55__R2_INV_1 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y55__R3_BUF_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y56__R0_BUF_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R0_INV_0 (.A(tie_lo_T12Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y56__R1_BUF_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R1_INV_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R2_INV_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y56__R2_INV_1 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y56__R3_BUF_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y57__R0_BUF_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R0_INV_0 (.A(tie_lo_T12Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y57__R1_BUF_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R1_INV_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R2_INV_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y57__R2_INV_1 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y57__R3_BUF_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y58__R0_BUF_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R0_INV_0 (.A(tie_lo_T12Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y58__R1_BUF_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R1_INV_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R2_INV_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y58__R2_INV_1 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y58__R3_BUF_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y59__R0_BUF_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R0_INV_0 (.A(tie_lo_T12Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y59__R1_BUF_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R1_INV_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R2_INV_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y59__R2_INV_1 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y59__R3_BUF_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y5__R0_BUF_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R0_INV_0 (.A(tie_lo_T12Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y5__R1_BUF_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R1_INV_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R2_INV_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y5__R2_INV_1 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y5__R3_BUF_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y60__R0_BUF_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R0_INV_0 (.A(tie_lo_T12Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y60__R1_BUF_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R1_INV_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R2_INV_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y60__R2_INV_1 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y60__R3_BUF_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y61__R0_BUF_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R0_INV_0 (.A(tie_lo_T12Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y61__R1_BUF_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R1_INV_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R2_INV_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y61__R2_INV_1 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y61__R3_BUF_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y62__R0_BUF_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R0_INV_0 (.A(tie_lo_T12Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y62__R1_BUF_0 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R1_INV_0 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R2_INV_0 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y62__R2_INV_1 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y62__R3_BUF_0 (.A(tie_lo_T12Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y63__R0_BUF_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R0_INV_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y63__R1_BUF_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R1_INV_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R2_INV_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y63__R2_INV_1 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y63__R3_BUF_0 (.A(tie_lo_T12Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y64__R0_BUF_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R0_INV_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y64__R1_BUF_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R1_INV_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R2_INV_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y64__R2_INV_1 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y64__R3_BUF_0 (.A(tie_lo_T12Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y65__R0_BUF_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R0_INV_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y65__R1_BUF_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R1_INV_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R2_INV_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y65__R2_INV_1 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y65__R3_BUF_0 (.A(tie_lo_T12Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y66__R0_BUF_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R0_INV_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y66__R1_BUF_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R1_INV_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R2_INV_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y66__R2_INV_1 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y66__R3_BUF_0 (.A(tie_lo_T12Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y67__R0_BUF_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R0_INV_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y67__R1_BUF_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R1_INV_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R2_INV_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y67__R2_INV_1 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y67__R3_BUF_0 (.A(tie_lo_T12Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y68__R0_BUF_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R0_INV_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y68__R1_BUF_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R1_INV_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R2_INV_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y68__R2_INV_1 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y68__R3_BUF_0 (.A(tie_lo_T12Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y69__R0_BUF_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R0_INV_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y69__R1_BUF_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R1_INV_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R2_INV_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y69__R2_INV_1 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y69__R3_BUF_0 (.A(tie_lo_T12Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y6__R0_BUF_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R0_INV_0 (.A(tie_lo_T12Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y6__R1_BUF_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R1_INV_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R2_INV_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y6__R2_INV_1 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y6__R3_BUF_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y70__R0_BUF_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R0_INV_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y70__R1_BUF_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R1_INV_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R2_INV_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y70__R2_INV_1 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y70__R3_BUF_0 (.A(tie_lo_T12Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y71__R0_BUF_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R0_INV_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y71__R1_BUF_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R1_INV_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R2_INV_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y71__R2_INV_1 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y71__R3_BUF_0 (.A(tie_lo_T12Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y72__R0_BUF_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R0_INV_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y72__R1_BUF_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R1_INV_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R2_INV_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y72__R2_INV_1 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y72__R3_BUF_0 (.A(tie_lo_T12Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y73__R0_BUF_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R0_INV_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y73__R1_BUF_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R1_INV_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R2_INV_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y73__R2_INV_1 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y73__R3_BUF_0 (.A(tie_lo_T12Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y74__R0_BUF_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R0_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y74__R1_BUF_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R1_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R2_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y74__R2_INV_1 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y74__R3_BUF_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y75__R0_BUF_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R0_INV_0 (.A(tie_lo_T12Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y75__R1_BUF_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R1_INV_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R2_INV_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y75__R2_INV_1 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y75__R3_BUF_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y76__R0_BUF_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R0_INV_0 (.A(tie_lo_T12Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y76__R1_BUF_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R1_INV_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R2_INV_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y76__R2_INV_1 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y76__R3_BUF_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y77__R0_BUF_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R0_INV_0 (.A(tie_lo_T12Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y77__R1_BUF_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R1_INV_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R2_INV_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y77__R2_INV_1 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y77__R3_BUF_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y78__R0_BUF_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R0_INV_0 (.A(tie_lo_T12Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y78__R1_BUF_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R1_INV_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R2_INV_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y78__R2_INV_1 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y78__R3_BUF_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y79__R0_BUF_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R0_INV_0 (.A(tie_lo_T12Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y79__R1_BUF_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R1_INV_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R2_INV_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y79__R2_INV_1 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y79__R3_BUF_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y7__R0_BUF_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R0_INV_0 (.A(tie_lo_T12Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y7__R1_BUF_0 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R1_INV_0 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R2_INV_0 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y7__R2_INV_1 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y7__R3_BUF_0 (.A(tie_lo_T12Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y80__R0_BUF_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R0_INV_0 (.A(tie_lo_T12Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y80__R1_BUF_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R1_INV_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R2_INV_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y80__R2_INV_1 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y80__R3_BUF_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y81__R0_BUF_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R0_INV_0 (.A(tie_lo_T12Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y81__R1_BUF_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R1_INV_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R2_INV_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y81__R2_INV_1 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y81__R3_BUF_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y82__R0_BUF_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R0_INV_0 (.A(tie_lo_T12Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y82__R1_BUF_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R1_INV_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R2_INV_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y82__R2_INV_1 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y82__R3_BUF_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y83__R0_BUF_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R0_INV_0 (.A(tie_lo_T12Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y83__R1_BUF_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R1_INV_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R2_INV_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y83__R2_INV_1 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y83__R3_BUF_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y84__R0_BUF_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R0_INV_0 (.A(tie_lo_T12Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y84__R1_BUF_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R1_INV_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R2_INV_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y84__R2_INV_1 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y84__R3_BUF_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y85__R0_BUF_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R0_INV_0 (.A(tie_lo_T12Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y85__R1_BUF_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R1_INV_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R2_INV_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y85__R2_INV_1 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y85__R3_BUF_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y86__R0_BUF_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R0_INV_0 (.A(tie_lo_T12Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y86__R1_BUF_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R1_INV_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R2_INV_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y86__R2_INV_1 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y86__R3_BUF_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y87__R0_BUF_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R0_INV_0 (.A(tie_lo_T12Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y87__R1_BUF_0 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R1_INV_0 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R2_INV_0 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y87__R2_INV_1 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y87__R3_BUF_0 (.A(tie_lo_T12Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y88__R0_BUF_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R0_INV_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y88__R1_BUF_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R1_INV_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R2_INV_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y88__R2_INV_1 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y88__R3_BUF_0 (.A(tie_lo_T12Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y89__R0_BUF_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R0_INV_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y89__R1_BUF_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R1_INV_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R2_INV_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y89__R2_INV_1 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y89__R3_BUF_0 (.A(tie_lo_T12Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y8__R0_BUF_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R0_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y8__R1_BUF_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R1_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R2_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y8__R2_INV_1 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y8__R3_BUF_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y9__R0_BUF_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R0_INV_0 (.A(tie_lo_T12Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y9__R1_BUF_0 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R1_INV_0 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T12Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R2_INV_0 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T12Y9__R2_INV_1 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T12Y9__R3_BUF_0 (.A(tie_lo_T12Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y0__R0_BUF_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R0_INV_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y0__R1_BUF_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R1_INV_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R2_INV_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y0__R2_INV_1 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y0__R3_BUF_0 (.A(tie_lo_T13Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y10__R0_BUF_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R0_INV_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y10__R1_BUF_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R1_INV_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R2_INV_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y10__R2_INV_1 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y10__R3_BUF_0 (.A(tie_lo_T13Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y11__R0_BUF_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R0_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y11__R1_BUF_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R1_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R2_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y11__R2_INV_1 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y11__R3_BUF_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y12__R0_BUF_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R0_INV_0 (.A(tie_lo_T13Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y12__R1_BUF_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R1_INV_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R2_INV_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y12__R2_INV_1 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y12__R3_BUF_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y13__R0_BUF_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R0_INV_0 (.A(tie_lo_T13Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y13__R1_BUF_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R1_INV_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R2_INV_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y13__R2_INV_1 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y13__R3_BUF_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y14__R0_BUF_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R0_INV_0 (.A(tie_lo_T13Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y14__R1_BUF_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R1_INV_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R2_INV_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y14__R2_INV_1 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y14__R3_BUF_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y15__R0_BUF_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R0_INV_0 (.A(tie_lo_T13Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y15__R1_BUF_0 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R1_INV_0 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R2_INV_0 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y15__R2_INV_1 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y15__R3_BUF_0 (.A(tie_lo_T13Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y16__R0_BUF_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R0_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y16__R1_BUF_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R1_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R2_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y16__R2_INV_1 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y16__R3_BUF_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y17__R0_BUF_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R0_INV_0 (.A(tie_lo_T13Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y17__R1_BUF_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R1_INV_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R2_INV_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y17__R2_INV_1 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y17__R3_BUF_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y18__R0_BUF_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R0_INV_0 (.A(tie_lo_T13Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y18__R1_BUF_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R1_INV_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R2_INV_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y18__R2_INV_1 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y18__R3_BUF_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y19__R0_BUF_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R0_INV_0 (.A(tie_lo_T13Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y19__R1_BUF_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R1_INV_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R2_INV_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y19__R2_INV_1 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y19__R3_BUF_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y1__R0_BUF_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R0_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y1__R1_BUF_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R1_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R2_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y1__R2_INV_1 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y1__R3_BUF_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y20__R0_BUF_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R0_INV_0 (.A(tie_lo_T13Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y20__R1_BUF_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R1_INV_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R2_INV_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y20__R2_INV_1 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y20__R3_BUF_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y21__R0_BUF_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R0_INV_0 (.A(tie_lo_T13Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y21__R1_BUF_0 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R1_INV_0 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R2_INV_0 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y21__R2_INV_1 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y21__R3_BUF_0 (.A(tie_lo_T13Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y22__R0_BUF_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R0_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y22__R1_BUF_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R1_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R2_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y22__R2_INV_1 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y22__R3_BUF_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y23__R0_BUF_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R0_INV_0 (.A(tie_lo_T13Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y23__R1_BUF_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R1_INV_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R2_INV_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y23__R2_INV_1 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y23__R3_BUF_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y24__R0_BUF_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R0_INV_0 (.A(tie_lo_T13Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y24__R1_BUF_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R1_INV_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R2_INV_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y24__R2_INV_1 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y24__R3_BUF_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y25__R0_BUF_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R0_INV_0 (.A(tie_lo_T13Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y25__R1_BUF_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R1_INV_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R2_INV_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y25__R2_INV_1 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y25__R3_BUF_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y26__R0_BUF_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R0_INV_0 (.A(tie_lo_T13Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y26__R1_BUF_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R1_INV_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R2_INV_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y26__R2_INV_1 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y26__R3_BUF_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y27__R0_BUF_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R0_INV_0 (.A(tie_lo_T13Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y27__R1_BUF_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R1_INV_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R2_INV_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y27__R2_INV_1 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y27__R3_BUF_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y28__R0_BUF_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R0_INV_0 (.A(tie_lo_T13Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y28__R1_BUF_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R1_INV_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R2_INV_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y28__R2_INV_1 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y28__R3_BUF_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y29__R0_BUF_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R0_INV_0 (.A(tie_lo_T13Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y29__R1_BUF_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R1_INV_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R2_INV_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y29__R2_INV_1 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y29__R3_BUF_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y2__R0_BUF_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R0_INV_0 (.A(tie_lo_T13Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y2__R1_BUF_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R1_INV_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R2_INV_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y2__R2_INV_1 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y2__R3_BUF_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y30__R0_BUF_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R0_INV_0 (.A(tie_lo_T13Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y30__R1_BUF_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R1_INV_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R2_INV_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y30__R2_INV_1 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y30__R3_BUF_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y31__R0_BUF_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R0_INV_0 (.A(tie_lo_T13Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y31__R1_BUF_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R1_INV_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R2_INV_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y31__R2_INV_1 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y31__R3_BUF_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y32__R0_BUF_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R0_INV_0 (.A(tie_lo_T13Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y32__R1_BUF_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R1_INV_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R2_INV_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y32__R2_INV_1 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y32__R3_BUF_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y33__R0_BUF_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R0_INV_0 (.A(tie_lo_T13Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y33__R1_BUF_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R1_INV_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R2_INV_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y33__R2_INV_1 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y33__R3_BUF_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y34__R0_BUF_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R0_INV_0 (.A(tie_lo_T13Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y34__R1_BUF_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R1_INV_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R2_INV_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y34__R2_INV_1 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y34__R3_BUF_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y35__R0_BUF_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R0_INV_0 (.A(tie_lo_T13Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y35__R1_BUF_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R1_INV_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R2_INV_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y35__R2_INV_1 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y35__R3_BUF_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y36__R0_BUF_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R0_INV_0 (.A(tie_lo_T13Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y36__R1_BUF_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R1_INV_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R2_INV_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y36__R2_INV_1 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y36__R3_BUF_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y37__R0_BUF_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R0_INV_0 (.A(tie_lo_T13Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y37__R1_BUF_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R1_INV_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R2_INV_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y37__R2_INV_1 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y37__R3_BUF_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y38__R0_BUF_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R0_INV_0 (.A(tie_lo_T13Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y38__R1_BUF_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R1_INV_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R2_INV_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y38__R2_INV_1 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y38__R3_BUF_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y39__R0_BUF_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R0_INV_0 (.A(tie_lo_T13Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y39__R1_BUF_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R1_INV_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R2_INV_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y39__R2_INV_1 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y39__R3_BUF_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y3__R0_BUF_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R0_INV_0 (.A(tie_lo_T13Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y3__R1_BUF_0 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R1_INV_0 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R2_INV_0 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y3__R2_INV_1 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y3__R3_BUF_0 (.A(tie_lo_T13Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y40__R0_BUF_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R0_INV_0 (.A(tie_lo_T13Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y40__R1_BUF_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R1_INV_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R2_INV_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y40__R2_INV_1 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y40__R3_BUF_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y41__R0_BUF_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R0_INV_0 (.A(tie_lo_T13Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y41__R1_BUF_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R1_INV_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R2_INV_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y41__R2_INV_1 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y41__R3_BUF_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y42__R0_BUF_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R0_INV_0 (.A(tie_lo_T13Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y42__R1_BUF_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R1_INV_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R2_INV_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y42__R2_INV_1 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y42__R3_BUF_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y43__R0_BUF_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R0_INV_0 (.A(tie_lo_T13Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y43__R1_BUF_0 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R1_INV_0 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R2_INV_0 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y43__R2_INV_1 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y43__R3_BUF_0 (.A(tie_lo_T13Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y44__R0_BUF_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R0_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y44__R1_BUF_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R1_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R2_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y44__R2_INV_1 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y44__R3_BUF_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y45__R0_BUF_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R0_INV_0 (.A(tie_lo_T13Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y45__R1_BUF_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R1_INV_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R2_INV_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y45__R2_INV_1 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y45__R3_BUF_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y46__R0_BUF_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R0_INV_0 (.A(tie_lo_T13Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y46__R1_BUF_0 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R1_INV_0 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R2_INV_0 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y46__R2_INV_1 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y46__R3_BUF_0 (.A(tie_lo_T13Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y47__R0_BUF_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R0_INV_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y47__R1_BUF_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R1_INV_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R2_INV_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y47__R2_INV_1 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y47__R3_BUF_0 (.A(tie_lo_T13Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y48__R0_BUF_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R0_INV_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y48__R1_BUF_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R1_INV_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R2_INV_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y48__R2_INV_1 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y48__R3_BUF_0 (.A(tie_lo_T13Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y49__R0_BUF_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R0_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y49__R1_BUF_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R1_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R2_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y49__R2_INV_1 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y49__R3_BUF_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y4__R0_BUF_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R0_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y4__R1_BUF_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R1_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R2_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y4__R2_INV_1 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y4__R3_BUF_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y50__R0_BUF_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R0_INV_0 (.A(tie_lo_T13Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y50__R1_BUF_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R1_INV_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R2_INV_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y50__R2_INV_1 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y50__R3_BUF_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y51__R0_BUF_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R0_INV_0 (.A(tie_lo_T13Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y51__R1_BUF_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R1_INV_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R2_INV_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y51__R2_INV_1 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y51__R3_BUF_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y52__R0_BUF_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R0_INV_0 (.A(tie_lo_T13Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y52__R1_BUF_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R1_INV_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R2_INV_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y52__R2_INV_1 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y52__R3_BUF_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y53__R0_BUF_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R0_INV_0 (.A(tie_lo_T13Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y53__R1_BUF_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R1_INV_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R2_INV_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y53__R2_INV_1 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y53__R3_BUF_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y54__R0_BUF_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R0_INV_0 (.A(tie_lo_T13Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y54__R1_BUF_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R1_INV_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R2_INV_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y54__R2_INV_1 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y54__R3_BUF_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y55__R0_BUF_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R0_INV_0 (.A(tie_lo_T13Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y55__R1_BUF_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R1_INV_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R2_INV_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y55__R2_INV_1 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y55__R3_BUF_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y56__R0_BUF_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R0_INV_0 (.A(tie_lo_T13Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y56__R1_BUF_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R1_INV_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R2_INV_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y56__R2_INV_1 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y56__R3_BUF_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y57__R0_BUF_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R0_INV_0 (.A(tie_lo_T13Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y57__R1_BUF_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R1_INV_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R2_INV_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y57__R2_INV_1 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y57__R3_BUF_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y58__R0_BUF_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R0_INV_0 (.A(tie_lo_T13Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y58__R1_BUF_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R1_INV_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R2_INV_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y58__R2_INV_1 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y58__R3_BUF_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y59__R0_BUF_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R0_INV_0 (.A(tie_lo_T13Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y59__R1_BUF_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R1_INV_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R2_INV_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y59__R2_INV_1 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y59__R3_BUF_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y5__R0_BUF_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R0_INV_0 (.A(tie_lo_T13Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y5__R1_BUF_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R1_INV_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R2_INV_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y5__R2_INV_1 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y5__R3_BUF_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y60__R0_BUF_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R0_INV_0 (.A(tie_lo_T13Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y60__R1_BUF_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R1_INV_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R2_INV_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y60__R2_INV_1 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y60__R3_BUF_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y61__R0_BUF_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R0_INV_0 (.A(tie_lo_T13Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y61__R1_BUF_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R1_INV_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R2_INV_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y61__R2_INV_1 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y61__R3_BUF_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y62__R0_BUF_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R0_INV_0 (.A(tie_lo_T13Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y62__R1_BUF_0 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R1_INV_0 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R2_INV_0 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y62__R2_INV_1 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y62__R3_BUF_0 (.A(tie_lo_T13Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y63__R0_BUF_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R0_INV_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y63__R1_BUF_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R1_INV_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R2_INV_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y63__R2_INV_1 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y63__R3_BUF_0 (.A(tie_lo_T13Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y64__R0_BUF_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R0_INV_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y64__R1_BUF_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R1_INV_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R2_INV_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y64__R2_INV_1 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y64__R3_BUF_0 (.A(tie_lo_T13Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y65__R0_BUF_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R0_INV_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y65__R1_BUF_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R1_INV_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R2_INV_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y65__R2_INV_1 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y65__R3_BUF_0 (.A(tie_lo_T13Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y66__R0_BUF_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R0_INV_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y66__R1_BUF_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R1_INV_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R2_INV_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y66__R2_INV_1 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y66__R3_BUF_0 (.A(tie_lo_T13Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y67__R0_BUF_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R0_INV_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y67__R1_BUF_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R1_INV_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R2_INV_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y67__R2_INV_1 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y67__R3_BUF_0 (.A(tie_lo_T13Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y68__R0_BUF_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R0_INV_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y68__R1_BUF_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R1_INV_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R2_INV_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y68__R2_INV_1 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y68__R3_BUF_0 (.A(tie_lo_T13Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y69__R0_BUF_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R0_INV_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y69__R1_BUF_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R1_INV_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R2_INV_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y69__R2_INV_1 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y69__R3_BUF_0 (.A(tie_lo_T13Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y6__R0_BUF_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R0_INV_0 (.A(tie_lo_T13Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y6__R1_BUF_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R1_INV_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R2_INV_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y6__R2_INV_1 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y6__R3_BUF_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y70__R0_BUF_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R0_INV_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y70__R1_BUF_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R1_INV_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R2_INV_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y70__R2_INV_1 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y70__R3_BUF_0 (.A(tie_lo_T13Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y71__R0_BUF_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R0_INV_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y71__R1_BUF_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R1_INV_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R2_INV_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y71__R2_INV_1 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y71__R3_BUF_0 (.A(tie_lo_T13Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y72__R0_BUF_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R0_INV_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y72__R1_BUF_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R1_INV_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R2_INV_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y72__R2_INV_1 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y72__R3_BUF_0 (.A(tie_lo_T13Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y73__R0_BUF_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R0_INV_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y73__R1_BUF_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R1_INV_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R2_INV_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y73__R2_INV_1 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y73__R3_BUF_0 (.A(tie_lo_T13Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y74__R0_BUF_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R0_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y74__R1_BUF_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R1_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R2_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y74__R2_INV_1 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y74__R3_BUF_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y75__R0_BUF_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R0_INV_0 (.A(tie_lo_T13Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y75__R1_BUF_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R1_INV_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R2_INV_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y75__R2_INV_1 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y75__R3_BUF_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y76__R0_BUF_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R0_INV_0 (.A(tie_lo_T13Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y76__R1_BUF_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R1_INV_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R2_INV_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y76__R2_INV_1 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y76__R3_BUF_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y77__R0_BUF_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R0_INV_0 (.A(tie_lo_T13Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y77__R1_BUF_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R1_INV_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R2_INV_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y77__R2_INV_1 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y77__R3_BUF_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y78__R0_BUF_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R0_INV_0 (.A(tie_lo_T13Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y78__R1_BUF_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R1_INV_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R2_INV_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y78__R2_INV_1 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y78__R3_BUF_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y79__R0_BUF_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R0_INV_0 (.A(tie_lo_T13Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y79__R1_BUF_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R1_INV_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R2_INV_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y79__R2_INV_1 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y79__R3_BUF_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y7__R0_BUF_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R0_INV_0 (.A(tie_lo_T13Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y7__R1_BUF_0 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R1_INV_0 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R2_INV_0 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y7__R2_INV_1 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y7__R3_BUF_0 (.A(tie_lo_T13Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y80__R0_BUF_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R0_INV_0 (.A(tie_lo_T13Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y80__R1_BUF_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R1_INV_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R2_INV_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y80__R2_INV_1 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y80__R3_BUF_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y81__R0_BUF_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R0_INV_0 (.A(tie_lo_T13Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y81__R1_BUF_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R1_INV_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R2_INV_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y81__R2_INV_1 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y81__R3_BUF_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y82__R0_BUF_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R0_INV_0 (.A(tie_lo_T13Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y82__R1_BUF_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R1_INV_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R2_INV_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y82__R2_INV_1 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y82__R3_BUF_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y83__R0_BUF_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R0_INV_0 (.A(tie_lo_T13Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y83__R1_BUF_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R1_INV_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R2_INV_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y83__R2_INV_1 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y83__R3_BUF_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y84__R0_BUF_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R0_INV_0 (.A(tie_lo_T13Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y84__R1_BUF_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R1_INV_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R2_INV_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y84__R2_INV_1 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y84__R3_BUF_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y85__R0_BUF_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R0_INV_0 (.A(tie_lo_T13Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y85__R1_BUF_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R1_INV_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R2_INV_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y85__R2_INV_1 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y85__R3_BUF_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y86__R0_BUF_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R0_INV_0 (.A(tie_lo_T13Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y86__R1_BUF_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R1_INV_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R2_INV_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y86__R2_INV_1 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y86__R3_BUF_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y87__R0_BUF_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R0_INV_0 (.A(tie_lo_T13Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y87__R1_BUF_0 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R1_INV_0 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R2_INV_0 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y87__R2_INV_1 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y87__R3_BUF_0 (.A(tie_lo_T13Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y88__R0_BUF_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R0_INV_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y88__R1_BUF_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R1_INV_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R2_INV_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y88__R2_INV_1 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y88__R3_BUF_0 (.A(tie_lo_T13Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y89__R0_BUF_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R0_INV_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y89__R1_BUF_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R1_INV_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R2_INV_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y89__R2_INV_1 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y89__R3_BUF_0 (.A(tie_lo_T13Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y8__R0_BUF_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R0_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y8__R1_BUF_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R1_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R2_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y8__R2_INV_1 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y8__R3_BUF_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y9__R0_BUF_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R0_INV_0 (.A(tie_lo_T13Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y9__R1_BUF_0 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R1_INV_0 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T13Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R2_INV_0 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T13Y9__R2_INV_1 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T13Y9__R3_BUF_0 (.A(tie_lo_T13Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y0__R0_BUF_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R0_INV_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y0__R1_BUF_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R1_INV_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R2_INV_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y0__R2_INV_1 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y0__R3_BUF_0 (.A(tie_lo_T14Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y10__R0_BUF_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R0_INV_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y10__R1_BUF_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R1_INV_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R2_INV_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y10__R2_INV_1 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y10__R3_BUF_0 (.A(tie_lo_T14Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y11__R0_BUF_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R0_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y11__R1_BUF_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R1_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R2_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y11__R2_INV_1 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y11__R3_BUF_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y12__R0_BUF_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R0_INV_0 (.A(tie_lo_T14Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y12__R1_BUF_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R1_INV_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R2_INV_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y12__R2_INV_1 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y12__R3_BUF_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y13__R0_BUF_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R0_INV_0 (.A(tie_lo_T14Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y13__R1_BUF_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R1_INV_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R2_INV_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y13__R2_INV_1 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y13__R3_BUF_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y14__R0_BUF_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R0_INV_0 (.A(tie_lo_T14Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y14__R1_BUF_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R1_INV_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R2_INV_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y14__R2_INV_1 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y14__R3_BUF_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y15__R0_BUF_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R0_INV_0 (.A(tie_lo_T14Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y15__R1_BUF_0 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R1_INV_0 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R2_INV_0 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y15__R2_INV_1 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y15__R3_BUF_0 (.A(tie_lo_T14Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y16__R0_BUF_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R0_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y16__R1_BUF_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R1_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R2_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y16__R2_INV_1 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y16__R3_BUF_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y17__R0_BUF_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R0_INV_0 (.A(tie_lo_T14Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y17__R1_BUF_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R1_INV_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R2_INV_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y17__R2_INV_1 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y17__R3_BUF_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y18__R0_BUF_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R0_INV_0 (.A(tie_lo_T14Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y18__R1_BUF_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R1_INV_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R2_INV_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y18__R2_INV_1 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y18__R3_BUF_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y19__R0_BUF_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R0_INV_0 (.A(tie_lo_T14Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y19__R1_BUF_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R1_INV_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R2_INV_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y19__R2_INV_1 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y19__R3_BUF_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y1__R0_BUF_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R0_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y1__R1_BUF_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R1_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R2_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y1__R2_INV_1 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y1__R3_BUF_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y20__R0_BUF_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R0_INV_0 (.A(tie_lo_T14Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y20__R1_BUF_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R1_INV_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R2_INV_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y20__R2_INV_1 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y20__R3_BUF_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y21__R0_BUF_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R0_INV_0 (.A(tie_lo_T14Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y21__R1_BUF_0 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R1_INV_0 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R2_INV_0 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y21__R2_INV_1 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y21__R3_BUF_0 (.A(tie_lo_T14Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y22__R0_BUF_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R0_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y22__R1_BUF_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R1_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R2_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y22__R2_INV_1 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y22__R3_BUF_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y23__R0_BUF_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R0_INV_0 (.A(tie_lo_T14Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y23__R1_BUF_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R1_INV_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R2_INV_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y23__R2_INV_1 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y23__R3_BUF_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y24__R0_BUF_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R0_INV_0 (.A(tie_lo_T14Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y24__R1_BUF_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R1_INV_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R2_INV_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y24__R2_INV_1 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y24__R3_BUF_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y25__R0_BUF_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R0_INV_0 (.A(tie_lo_T14Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y25__R1_BUF_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R1_INV_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R2_INV_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y25__R2_INV_1 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y25__R3_BUF_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y26__R0_BUF_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R0_INV_0 (.A(tie_lo_T14Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y26__R1_BUF_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R1_INV_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R2_INV_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y26__R2_INV_1 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y26__R3_BUF_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y27__R0_BUF_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R0_INV_0 (.A(tie_lo_T14Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y27__R1_BUF_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R1_INV_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R2_INV_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y27__R2_INV_1 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y27__R3_BUF_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y28__R0_BUF_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R0_INV_0 (.A(tie_lo_T14Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y28__R1_BUF_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R1_INV_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R2_INV_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y28__R2_INV_1 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y28__R3_BUF_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y29__R0_BUF_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R0_INV_0 (.A(tie_lo_T14Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y29__R1_BUF_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R1_INV_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R2_INV_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y29__R2_INV_1 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y29__R3_BUF_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y2__R0_BUF_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R0_INV_0 (.A(tie_lo_T14Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y2__R1_BUF_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R1_INV_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R2_INV_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y2__R2_INV_1 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y2__R3_BUF_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y30__R0_BUF_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R0_INV_0 (.A(tie_lo_T14Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y30__R1_BUF_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R1_INV_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R2_INV_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y30__R2_INV_1 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y30__R3_BUF_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y31__R0_BUF_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R0_INV_0 (.A(tie_lo_T14Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y31__R1_BUF_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R1_INV_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R2_INV_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y31__R2_INV_1 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y31__R3_BUF_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y32__R0_BUF_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R0_INV_0 (.A(tie_lo_T14Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y32__R1_BUF_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R1_INV_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R2_INV_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y32__R2_INV_1 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y32__R3_BUF_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y33__R0_BUF_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R0_INV_0 (.A(tie_lo_T14Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y33__R1_BUF_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R1_INV_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R2_INV_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y33__R2_INV_1 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y33__R3_BUF_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y34__R0_BUF_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R0_INV_0 (.A(tie_lo_T14Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y34__R1_BUF_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R1_INV_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R2_INV_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y34__R2_INV_1 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y34__R3_BUF_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y35__R0_BUF_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R0_INV_0 (.A(tie_lo_T14Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y35__R1_BUF_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R1_INV_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R2_INV_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y35__R2_INV_1 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y35__R3_BUF_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y36__R0_BUF_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R0_INV_0 (.A(tie_lo_T14Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y36__R1_BUF_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R1_INV_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R2_INV_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y36__R2_INV_1 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y36__R3_BUF_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y37__R0_BUF_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R0_INV_0 (.A(tie_lo_T14Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y37__R1_BUF_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R1_INV_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R2_INV_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y37__R2_INV_1 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y37__R3_BUF_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y38__R0_BUF_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R0_INV_0 (.A(tie_lo_T14Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y38__R1_BUF_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R1_INV_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R2_INV_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y38__R2_INV_1 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y38__R3_BUF_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y39__R0_BUF_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R0_INV_0 (.A(tie_lo_T14Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y39__R1_BUF_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R1_INV_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R2_INV_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y39__R2_INV_1 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y39__R3_BUF_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y3__R0_BUF_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R0_INV_0 (.A(tie_lo_T14Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y3__R1_BUF_0 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R1_INV_0 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R2_INV_0 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y3__R2_INV_1 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y3__R3_BUF_0 (.A(tie_lo_T14Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y40__R0_BUF_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R0_INV_0 (.A(tie_lo_T14Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y40__R1_BUF_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R1_INV_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R2_INV_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y40__R2_INV_1 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y40__R3_BUF_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y41__R0_BUF_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R0_INV_0 (.A(tie_lo_T14Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y41__R1_BUF_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R1_INV_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R2_INV_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y41__R2_INV_1 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y41__R3_BUF_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y42__R0_BUF_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R0_INV_0 (.A(tie_lo_T14Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y42__R1_BUF_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R1_INV_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R2_INV_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y42__R2_INV_1 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y42__R3_BUF_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y43__R0_BUF_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R0_INV_0 (.A(tie_lo_T14Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y43__R1_BUF_0 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R1_INV_0 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R2_INV_0 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y43__R2_INV_1 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y43__R3_BUF_0 (.A(tie_lo_T14Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y44__R0_BUF_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R0_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y44__R1_BUF_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R1_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R2_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y44__R2_INV_1 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y44__R3_BUF_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y45__R0_BUF_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R0_INV_0 (.A(tie_lo_T14Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y45__R1_BUF_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R1_INV_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R2_INV_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y45__R2_INV_1 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y45__R3_BUF_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y46__R0_BUF_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R0_INV_0 (.A(tie_lo_T14Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y46__R1_BUF_0 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R1_INV_0 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R2_INV_0 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y46__R2_INV_1 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y46__R3_BUF_0 (.A(tie_lo_T14Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y47__R0_BUF_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R0_INV_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y47__R1_BUF_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R1_INV_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R2_INV_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y47__R2_INV_1 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y47__R3_BUF_0 (.A(tie_lo_T14Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y48__R0_BUF_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R0_INV_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y48__R1_BUF_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R1_INV_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R2_INV_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y48__R2_INV_1 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y48__R3_BUF_0 (.A(tie_lo_T14Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y49__R0_BUF_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R0_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y49__R1_BUF_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R1_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R2_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y49__R2_INV_1 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y49__R3_BUF_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y4__R0_BUF_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R0_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y4__R1_BUF_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R1_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R2_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y4__R2_INV_1 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y4__R3_BUF_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y50__R0_BUF_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R0_INV_0 (.A(tie_lo_T14Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y50__R1_BUF_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R1_INV_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R2_INV_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y50__R2_INV_1 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y50__R3_BUF_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y51__R0_BUF_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R0_INV_0 (.A(tie_lo_T14Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y51__R1_BUF_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R1_INV_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R2_INV_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y51__R2_INV_1 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y51__R3_BUF_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y52__R0_BUF_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R0_INV_0 (.A(tie_lo_T14Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y52__R1_BUF_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R1_INV_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R2_INV_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y52__R2_INV_1 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y52__R3_BUF_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y53__R0_BUF_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R0_INV_0 (.A(tie_lo_T14Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y53__R1_BUF_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R1_INV_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R2_INV_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y53__R2_INV_1 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y53__R3_BUF_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y54__R0_BUF_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R0_INV_0 (.A(tie_lo_T14Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y54__R1_BUF_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R1_INV_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R2_INV_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y54__R2_INV_1 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y54__R3_BUF_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y55__R0_BUF_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R0_INV_0 (.A(tie_lo_T14Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y55__R1_BUF_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R1_INV_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R2_INV_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y55__R2_INV_1 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y55__R3_BUF_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y56__R0_BUF_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R0_INV_0 (.A(tie_lo_T14Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y56__R1_BUF_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R1_INV_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R2_INV_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y56__R2_INV_1 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y56__R3_BUF_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y57__R0_BUF_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R0_INV_0 (.A(tie_lo_T14Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y57__R1_BUF_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R1_INV_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R2_INV_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y57__R2_INV_1 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y57__R3_BUF_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y58__R0_BUF_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R0_INV_0 (.A(tie_lo_T14Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y58__R1_BUF_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R1_INV_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R2_INV_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y58__R2_INV_1 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y58__R3_BUF_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y59__R0_BUF_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R0_INV_0 (.A(tie_lo_T14Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y59__R1_BUF_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R1_INV_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R2_INV_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y59__R2_INV_1 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y59__R3_BUF_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y5__R0_BUF_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R0_INV_0 (.A(tie_lo_T14Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y5__R1_BUF_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R1_INV_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R2_INV_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y5__R2_INV_1 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y5__R3_BUF_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y60__R0_BUF_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R0_INV_0 (.A(tie_lo_T14Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y60__R1_BUF_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R1_INV_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R2_INV_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y60__R2_INV_1 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y60__R3_BUF_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y61__R0_BUF_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R0_INV_0 (.A(tie_lo_T14Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y61__R1_BUF_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R1_INV_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R2_INV_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y61__R2_INV_1 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y61__R3_BUF_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y62__R0_BUF_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R0_INV_0 (.A(tie_lo_T14Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y62__R1_BUF_0 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R1_INV_0 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R2_INV_0 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y62__R2_INV_1 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y62__R3_BUF_0 (.A(tie_lo_T14Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y63__R0_BUF_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R0_INV_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y63__R1_BUF_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R1_INV_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R2_INV_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y63__R2_INV_1 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y63__R3_BUF_0 (.A(tie_lo_T14Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y64__R0_BUF_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R0_INV_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y64__R1_BUF_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R1_INV_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R2_INV_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y64__R2_INV_1 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y64__R3_BUF_0 (.A(tie_lo_T14Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y65__R0_BUF_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R0_INV_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y65__R1_BUF_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R1_INV_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R2_INV_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y65__R2_INV_1 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y65__R3_BUF_0 (.A(tie_lo_T14Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y66__R0_BUF_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R0_INV_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y66__R1_BUF_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R1_INV_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R2_INV_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y66__R2_INV_1 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y66__R3_BUF_0 (.A(tie_lo_T14Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y67__R0_BUF_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R0_INV_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y67__R1_BUF_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R1_INV_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R2_INV_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y67__R2_INV_1 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y67__R3_BUF_0 (.A(tie_lo_T14Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y68__R0_BUF_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R0_INV_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y68__R1_BUF_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R1_INV_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R2_INV_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y68__R2_INV_1 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y68__R3_BUF_0 (.A(tie_lo_T14Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y69__R0_BUF_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R0_INV_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y69__R1_BUF_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R1_INV_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R2_INV_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y69__R2_INV_1 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y69__R3_BUF_0 (.A(tie_lo_T14Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y6__R0_BUF_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R0_INV_0 (.A(tie_lo_T14Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y6__R1_BUF_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R1_INV_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R2_INV_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y6__R2_INV_1 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y6__R3_BUF_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y70__R0_BUF_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R0_INV_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y70__R1_BUF_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R1_INV_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R2_INV_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y70__R2_INV_1 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y70__R3_BUF_0 (.A(tie_lo_T14Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y71__R0_BUF_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R0_INV_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y71__R1_BUF_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R1_INV_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R2_INV_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y71__R2_INV_1 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y71__R3_BUF_0 (.A(tie_lo_T14Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y72__R0_BUF_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R0_INV_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y72__R1_BUF_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R1_INV_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R2_INV_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y72__R2_INV_1 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y72__R3_BUF_0 (.A(tie_lo_T14Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y73__R0_BUF_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R0_INV_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y73__R1_BUF_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R1_INV_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R2_INV_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y73__R2_INV_1 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y73__R3_BUF_0 (.A(tie_lo_T14Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y74__R0_BUF_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R0_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y74__R1_BUF_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R1_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R2_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y74__R2_INV_1 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y74__R3_BUF_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y75__R0_BUF_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R0_INV_0 (.A(tie_lo_T14Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y75__R1_BUF_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R1_INV_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R2_INV_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y75__R2_INV_1 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y75__R3_BUF_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y76__R0_BUF_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R0_INV_0 (.A(tie_lo_T14Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y76__R1_BUF_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R1_INV_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R2_INV_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y76__R2_INV_1 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y76__R3_BUF_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y77__R0_BUF_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R0_INV_0 (.A(tie_lo_T14Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y77__R1_BUF_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R1_INV_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R2_INV_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y77__R2_INV_1 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y77__R3_BUF_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y78__R0_BUF_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R0_INV_0 (.A(tie_lo_T14Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y78__R1_BUF_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R1_INV_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R2_INV_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y78__R2_INV_1 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y78__R3_BUF_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y79__R0_BUF_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R0_INV_0 (.A(tie_lo_T14Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y79__R1_BUF_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R1_INV_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R2_INV_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y79__R2_INV_1 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y79__R3_BUF_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y7__R0_BUF_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R0_INV_0 (.A(tie_lo_T14Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y7__R1_BUF_0 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R1_INV_0 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R2_INV_0 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y7__R2_INV_1 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y7__R3_BUF_0 (.A(tie_lo_T14Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y80__R0_BUF_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R0_INV_0 (.A(tie_lo_T14Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y80__R1_BUF_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R1_INV_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R2_INV_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y80__R2_INV_1 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y80__R3_BUF_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y81__R0_BUF_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R0_INV_0 (.A(tie_lo_T14Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y81__R1_BUF_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R1_INV_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R2_INV_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y81__R2_INV_1 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y81__R3_BUF_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y82__R0_BUF_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R0_INV_0 (.A(tie_lo_T14Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y82__R1_BUF_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R1_INV_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R2_INV_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y82__R2_INV_1 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y82__R3_BUF_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y83__R0_BUF_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R0_INV_0 (.A(tie_lo_T14Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y83__R1_BUF_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R1_INV_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R2_INV_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y83__R2_INV_1 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y83__R3_BUF_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y84__R0_BUF_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R0_INV_0 (.A(tie_lo_T14Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y84__R1_BUF_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R1_INV_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R2_INV_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y84__R2_INV_1 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y84__R3_BUF_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y85__R0_BUF_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R0_INV_0 (.A(tie_lo_T14Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y85__R1_BUF_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R1_INV_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R2_INV_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y85__R2_INV_1 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y85__R3_BUF_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y86__R0_BUF_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R0_INV_0 (.A(tie_lo_T14Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y86__R1_BUF_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R1_INV_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R2_INV_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y86__R2_INV_1 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y86__R3_BUF_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y87__R0_BUF_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R0_INV_0 (.A(tie_lo_T14Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y87__R1_BUF_0 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R1_INV_0 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R2_INV_0 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y87__R2_INV_1 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y87__R3_BUF_0 (.A(tie_lo_T14Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y88__R0_BUF_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R0_INV_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y88__R1_BUF_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R1_INV_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R2_INV_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y88__R2_INV_1 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y88__R3_BUF_0 (.A(tie_lo_T14Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y89__R0_BUF_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R0_INV_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y89__R1_BUF_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R1_INV_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R2_INV_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y89__R2_INV_1 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y89__R3_BUF_0 (.A(tie_lo_T14Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y8__R0_BUF_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R0_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y8__R1_BUF_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R1_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R2_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y8__R2_INV_1 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y8__R3_BUF_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y9__R0_BUF_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R0_INV_0 (.A(tie_lo_T14Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y9__R1_BUF_0 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R1_INV_0 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T14Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R2_INV_0 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T14Y9__R2_INV_1 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T14Y9__R3_BUF_0 (.A(tie_lo_T14Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y0__R0_BUF_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R0_INV_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y0__R1_BUF_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R1_INV_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R2_INV_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y0__R2_INV_1 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y0__R3_BUF_0 (.A(tie_lo_T15Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y10__R0_BUF_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R0_INV_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y10__R1_BUF_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R1_INV_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R2_INV_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y10__R2_INV_1 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y10__R3_BUF_0 (.A(tie_lo_T15Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y11__R0_BUF_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R0_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y11__R1_BUF_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R1_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R2_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y11__R2_INV_1 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y11__R3_BUF_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y12__R0_BUF_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R0_INV_0 (.A(tie_lo_T15Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y12__R1_BUF_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R1_INV_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R2_INV_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y12__R2_INV_1 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y12__R3_BUF_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y13__R0_BUF_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R0_INV_0 (.A(tie_lo_T15Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y13__R1_BUF_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R1_INV_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R2_INV_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y13__R2_INV_1 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y13__R3_BUF_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y14__R0_BUF_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R0_INV_0 (.A(tie_lo_T15Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y14__R1_BUF_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R1_INV_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R2_INV_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y14__R2_INV_1 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y14__R3_BUF_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y15__R0_BUF_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R0_INV_0 (.A(tie_lo_T15Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y15__R1_BUF_0 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R1_INV_0 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R2_INV_0 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y15__R2_INV_1 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y15__R3_BUF_0 (.A(tie_lo_T15Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y16__R0_BUF_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R0_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y16__R1_BUF_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R1_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R2_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y16__R2_INV_1 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y16__R3_BUF_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y17__R0_BUF_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R0_INV_0 (.A(tie_lo_T15Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y17__R1_BUF_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R1_INV_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R2_INV_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y17__R2_INV_1 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y17__R3_BUF_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y18__R0_BUF_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R0_INV_0 (.A(tie_lo_T15Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y18__R1_BUF_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R1_INV_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R2_INV_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y18__R2_INV_1 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y18__R3_BUF_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y19__R0_BUF_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R0_INV_0 (.A(tie_lo_T15Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y19__R1_BUF_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R1_INV_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R2_INV_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y19__R2_INV_1 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y19__R3_BUF_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y1__R0_BUF_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R0_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y1__R1_BUF_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R1_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R2_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y1__R2_INV_1 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y1__R3_BUF_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y20__R0_BUF_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R0_INV_0 (.A(tie_lo_T15Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y20__R1_BUF_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R1_INV_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R2_INV_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y20__R2_INV_1 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y20__R3_BUF_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y21__R0_BUF_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R0_INV_0 (.A(tie_lo_T15Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y21__R1_BUF_0 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R1_INV_0 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R2_INV_0 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y21__R2_INV_1 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y21__R3_BUF_0 (.A(tie_lo_T15Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y22__R0_BUF_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R0_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y22__R1_BUF_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R1_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R2_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y22__R2_INV_1 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y22__R3_BUF_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y23__R0_BUF_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R0_INV_0 (.A(tie_lo_T15Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y23__R1_BUF_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R1_INV_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R2_INV_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y23__R2_INV_1 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y23__R3_BUF_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y24__R0_BUF_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R0_INV_0 (.A(tie_lo_T15Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y24__R1_BUF_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R1_INV_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R2_INV_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y24__R2_INV_1 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y24__R3_BUF_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y25__R0_BUF_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R0_INV_0 (.A(tie_lo_T15Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y25__R1_BUF_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R1_INV_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R2_INV_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y25__R2_INV_1 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y25__R3_BUF_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y26__R0_BUF_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R0_INV_0 (.A(tie_lo_T15Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y26__R1_BUF_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R1_INV_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R2_INV_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y26__R2_INV_1 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y26__R3_BUF_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y27__R0_BUF_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R0_INV_0 (.A(tie_lo_T15Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y27__R1_BUF_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R1_INV_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R2_INV_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y27__R2_INV_1 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y27__R3_BUF_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y28__R0_BUF_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R0_INV_0 (.A(tie_lo_T15Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y28__R1_BUF_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R1_INV_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R2_INV_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y28__R2_INV_1 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y28__R3_BUF_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y29__R0_BUF_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R0_INV_0 (.A(tie_lo_T15Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y29__R1_BUF_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R1_INV_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R2_INV_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y29__R2_INV_1 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y29__R3_BUF_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y2__R0_BUF_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R0_INV_0 (.A(tie_lo_T15Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y2__R1_BUF_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R1_INV_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R2_INV_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y2__R2_INV_1 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y2__R3_BUF_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y30__R0_BUF_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R0_INV_0 (.A(tie_lo_T15Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y30__R1_BUF_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R1_INV_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R2_INV_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y30__R2_INV_1 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y30__R3_BUF_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y31__R0_BUF_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R0_INV_0 (.A(tie_lo_T15Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y31__R1_BUF_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R1_INV_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R2_INV_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y31__R2_INV_1 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y31__R3_BUF_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y32__R0_BUF_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R0_INV_0 (.A(tie_lo_T15Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y32__R1_BUF_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R1_INV_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R2_INV_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y32__R2_INV_1 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y32__R3_BUF_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y33__R0_BUF_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R0_INV_0 (.A(tie_lo_T15Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y33__R1_BUF_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R1_INV_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R2_INV_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y33__R2_INV_1 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y33__R3_BUF_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y34__R0_BUF_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R0_INV_0 (.A(tie_lo_T15Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y34__R1_BUF_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R1_INV_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R2_INV_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y34__R2_INV_1 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y34__R3_BUF_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y35__R0_BUF_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R0_INV_0 (.A(tie_lo_T15Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y35__R1_BUF_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R1_INV_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R2_INV_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y35__R2_INV_1 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y35__R3_BUF_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y36__R0_BUF_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R0_INV_0 (.A(tie_lo_T15Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y36__R1_BUF_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R1_INV_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R2_INV_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y36__R2_INV_1 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y36__R3_BUF_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y37__R0_BUF_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R0_INV_0 (.A(tie_lo_T15Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y37__R1_BUF_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R1_INV_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R2_INV_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y37__R2_INV_1 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y37__R3_BUF_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y38__R0_BUF_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R0_INV_0 (.A(tie_lo_T15Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y38__R1_BUF_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R1_INV_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R2_INV_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y38__R2_INV_1 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y38__R3_BUF_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y39__R0_BUF_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R0_INV_0 (.A(tie_lo_T15Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y39__R1_BUF_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R1_INV_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R2_INV_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y39__R2_INV_1 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y39__R3_BUF_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y3__R0_BUF_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R0_INV_0 (.A(tie_lo_T15Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y3__R1_BUF_0 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R1_INV_0 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R2_INV_0 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y3__R2_INV_1 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y3__R3_BUF_0 (.A(tie_lo_T15Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y40__R0_BUF_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R0_INV_0 (.A(tie_lo_T15Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y40__R1_BUF_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R1_INV_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R2_INV_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y40__R2_INV_1 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y40__R3_BUF_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y41__R0_BUF_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R0_INV_0 (.A(tie_lo_T15Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y41__R1_BUF_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R1_INV_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R2_INV_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y41__R2_INV_1 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y41__R3_BUF_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y42__R0_BUF_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R0_INV_0 (.A(tie_lo_T15Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y42__R1_BUF_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R1_INV_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R2_INV_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y42__R2_INV_1 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y42__R3_BUF_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y43__R0_BUF_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R0_INV_0 (.A(tie_lo_T15Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y43__R1_BUF_0 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R1_INV_0 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R2_INV_0 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y43__R2_INV_1 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y43__R3_BUF_0 (.A(tie_lo_T15Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y44__R0_BUF_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R0_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y44__R1_BUF_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R1_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R2_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y44__R2_INV_1 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y44__R3_BUF_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y45__R0_BUF_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R0_INV_0 (.A(tie_lo_T15Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y45__R1_BUF_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R1_INV_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R2_INV_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y45__R2_INV_1 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y45__R3_BUF_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y46__R0_BUF_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R0_INV_0 (.A(tie_lo_T15Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y46__R1_BUF_0 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R1_INV_0 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R2_INV_0 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y46__R2_INV_1 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y46__R3_BUF_0 (.A(tie_lo_T15Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y47__R0_BUF_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R0_INV_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y47__R1_BUF_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R1_INV_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R2_INV_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y47__R2_INV_1 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y47__R3_BUF_0 (.A(tie_lo_T15Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y48__R0_BUF_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R0_INV_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y48__R1_BUF_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R1_INV_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R2_INV_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y48__R2_INV_1 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y48__R3_BUF_0 (.A(tie_lo_T15Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y49__R0_BUF_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R0_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y49__R1_BUF_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R1_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R2_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y49__R2_INV_1 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y49__R3_BUF_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y4__R0_BUF_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R0_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y4__R1_BUF_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R1_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R2_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y4__R2_INV_1 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y4__R3_BUF_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y50__R0_BUF_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R0_INV_0 (.A(tie_lo_T15Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y50__R1_BUF_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R1_INV_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R2_INV_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y50__R2_INV_1 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y50__R3_BUF_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y51__R0_BUF_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R0_INV_0 (.A(tie_lo_T15Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y51__R1_BUF_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R1_INV_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R2_INV_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y51__R2_INV_1 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y51__R3_BUF_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y52__R0_BUF_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R0_INV_0 (.A(tie_lo_T15Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y52__R1_BUF_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R1_INV_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R2_INV_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y52__R2_INV_1 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y52__R3_BUF_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y53__R0_BUF_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R0_INV_0 (.A(tie_lo_T15Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y53__R1_BUF_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R1_INV_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R2_INV_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y53__R2_INV_1 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y53__R3_BUF_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y54__R0_BUF_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R0_INV_0 (.A(tie_lo_T15Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y54__R1_BUF_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R1_INV_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R2_INV_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y54__R2_INV_1 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y54__R3_BUF_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y55__R0_BUF_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R0_INV_0 (.A(tie_lo_T15Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y55__R1_BUF_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R1_INV_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R2_INV_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y55__R2_INV_1 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y55__R3_BUF_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y56__R0_BUF_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R0_INV_0 (.A(tie_lo_T15Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y56__R1_BUF_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R1_INV_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R2_INV_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y56__R2_INV_1 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y56__R3_BUF_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y57__R0_BUF_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R0_INV_0 (.A(tie_lo_T15Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y57__R1_BUF_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R1_INV_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R2_INV_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y57__R2_INV_1 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y57__R3_BUF_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y58__R0_BUF_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R0_INV_0 (.A(tie_lo_T15Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y58__R1_BUF_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R1_INV_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R2_INV_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y58__R2_INV_1 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y58__R3_BUF_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y59__R0_BUF_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R0_INV_0 (.A(tie_lo_T15Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y59__R1_BUF_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R1_INV_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R2_INV_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y59__R2_INV_1 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y59__R3_BUF_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y5__R0_BUF_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R0_INV_0 (.A(tie_lo_T15Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y5__R1_BUF_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R1_INV_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R2_INV_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y5__R2_INV_1 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y5__R3_BUF_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y60__R0_BUF_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R0_INV_0 (.A(tie_lo_T15Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y60__R1_BUF_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R1_INV_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R2_INV_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y60__R2_INV_1 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y60__R3_BUF_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y61__R0_BUF_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R0_INV_0 (.A(tie_lo_T15Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y61__R1_BUF_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R1_INV_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R2_INV_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y61__R2_INV_1 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y61__R3_BUF_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y62__R0_BUF_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R0_INV_0 (.A(tie_lo_T15Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y62__R1_BUF_0 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R1_INV_0 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R2_INV_0 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y62__R2_INV_1 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y62__R3_BUF_0 (.A(tie_lo_T15Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y63__R0_BUF_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R0_INV_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y63__R1_BUF_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R1_INV_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R2_INV_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y63__R2_INV_1 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y63__R3_BUF_0 (.A(tie_lo_T15Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y64__R0_BUF_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R0_INV_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y64__R1_BUF_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R1_INV_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R2_INV_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y64__R2_INV_1 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y64__R3_BUF_0 (.A(tie_lo_T15Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y65__R0_BUF_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R0_INV_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y65__R1_BUF_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R1_INV_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R2_INV_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y65__R2_INV_1 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y65__R3_BUF_0 (.A(tie_lo_T15Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y66__R0_BUF_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R0_INV_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y66__R1_BUF_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R1_INV_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R2_INV_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y66__R2_INV_1 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y66__R3_BUF_0 (.A(tie_lo_T15Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y67__R0_BUF_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R0_INV_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y67__R1_BUF_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R1_INV_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R2_INV_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y67__R2_INV_1 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y67__R3_BUF_0 (.A(tie_lo_T15Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y68__R0_BUF_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R0_INV_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y68__R1_BUF_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R1_INV_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R2_INV_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y68__R2_INV_1 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y68__R3_BUF_0 (.A(tie_lo_T15Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y69__R0_BUF_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R0_INV_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y69__R1_BUF_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R1_INV_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R2_INV_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y69__R2_INV_1 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y69__R3_BUF_0 (.A(tie_lo_T15Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y6__R0_BUF_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R0_INV_0 (.A(tie_lo_T15Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y6__R1_BUF_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R1_INV_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R2_INV_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y6__R2_INV_1 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y6__R3_BUF_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y70__R0_BUF_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R0_INV_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y70__R1_BUF_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R1_INV_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R2_INV_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y70__R2_INV_1 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y70__R3_BUF_0 (.A(tie_lo_T15Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y71__R0_BUF_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R0_INV_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y71__R1_BUF_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R1_INV_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R2_INV_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y71__R2_INV_1 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y71__R3_BUF_0 (.A(tie_lo_T15Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y72__R0_BUF_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R0_INV_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y72__R1_BUF_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R1_INV_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R2_INV_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y72__R2_INV_1 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y72__R3_BUF_0 (.A(tie_lo_T15Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y73__R0_BUF_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R0_INV_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y73__R1_BUF_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R1_INV_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R2_INV_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y73__R2_INV_1 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y73__R3_BUF_0 (.A(tie_lo_T15Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y74__R0_BUF_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R0_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y74__R1_BUF_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R1_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R2_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y74__R2_INV_1 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y74__R3_BUF_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y75__R0_BUF_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R0_INV_0 (.A(tie_lo_T15Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y75__R1_BUF_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R1_INV_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R2_INV_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y75__R2_INV_1 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y75__R3_BUF_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y76__R0_BUF_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R0_INV_0 (.A(tie_lo_T15Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y76__R1_BUF_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R1_INV_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R2_INV_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y76__R2_INV_1 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y76__R3_BUF_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y77__R0_BUF_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R0_INV_0 (.A(tie_lo_T15Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y77__R1_BUF_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R1_INV_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R2_INV_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y77__R2_INV_1 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y77__R3_BUF_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y78__R0_BUF_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R0_INV_0 (.A(tie_lo_T15Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y78__R1_BUF_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R1_INV_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R2_INV_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y78__R2_INV_1 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y78__R3_BUF_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y79__R0_BUF_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R0_INV_0 (.A(tie_lo_T15Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y79__R1_BUF_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R1_INV_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R2_INV_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y79__R2_INV_1 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y79__R3_BUF_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y7__R0_BUF_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R0_INV_0 (.A(tie_lo_T15Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y7__R1_BUF_0 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R1_INV_0 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R2_INV_0 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y7__R2_INV_1 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y7__R3_BUF_0 (.A(tie_lo_T15Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y80__R0_BUF_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R0_INV_0 (.A(tie_lo_T15Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y80__R1_BUF_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R1_INV_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R2_INV_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y80__R2_INV_1 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y80__R3_BUF_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y81__R0_BUF_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R0_INV_0 (.A(tie_lo_T15Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y81__R1_BUF_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R1_INV_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R2_INV_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y81__R2_INV_1 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y81__R3_BUF_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y82__R0_BUF_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R0_INV_0 (.A(tie_lo_T15Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y82__R1_BUF_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R1_INV_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R2_INV_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y82__R2_INV_1 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y82__R3_BUF_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y83__R0_BUF_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R0_INV_0 (.A(tie_lo_T15Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y83__R1_BUF_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R1_INV_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R2_INV_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y83__R2_INV_1 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y83__R3_BUF_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y84__R0_BUF_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R0_INV_0 (.A(tie_lo_T15Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y84__R1_BUF_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R1_INV_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R2_INV_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y84__R2_INV_1 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y84__R3_BUF_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y85__R0_BUF_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R0_INV_0 (.A(tie_lo_T15Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y85__R1_BUF_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R1_INV_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R2_INV_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y85__R2_INV_1 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y85__R3_BUF_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y86__R0_BUF_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R0_INV_0 (.A(tie_lo_T15Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y86__R1_BUF_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R1_INV_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R2_INV_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y86__R2_INV_1 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y86__R3_BUF_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y87__R0_BUF_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R0_INV_0 (.A(tie_lo_T15Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y87__R1_BUF_0 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R1_INV_0 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R2_INV_0 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y87__R2_INV_1 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y87__R3_BUF_0 (.A(tie_lo_T15Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y88__R0_BUF_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R0_INV_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y88__R1_BUF_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R1_INV_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R2_INV_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y88__R2_INV_1 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y88__R3_BUF_0 (.A(tie_lo_T15Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y89__R0_BUF_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R0_INV_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y89__R1_BUF_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R1_INV_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R2_INV_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y89__R2_INV_1 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y89__R3_BUF_0 (.A(tie_lo_T15Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y8__R0_BUF_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R0_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y8__R1_BUF_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R1_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R2_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y8__R2_INV_1 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y8__R3_BUF_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y9__R0_BUF_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R0_INV_0 (.A(tie_lo_T15Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y9__R1_BUF_0 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R1_INV_0 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T15Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R2_INV_0 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T15Y9__R2_INV_1 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T15Y9__R3_BUF_0 (.A(tie_lo_T15Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y0__R0_BUF_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R0_INV_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y0__R1_BUF_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R1_INV_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R2_INV_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y0__R2_INV_1 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y0__R3_BUF_0 (.A(tie_lo_T16Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y10__R0_BUF_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R0_INV_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y10__R1_BUF_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R1_INV_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R2_INV_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y10__R2_INV_1 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y10__R3_BUF_0 (.A(tie_lo_T16Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y11__R0_BUF_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R0_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y11__R1_BUF_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R1_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R2_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y11__R2_INV_1 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y11__R3_BUF_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y12__R0_BUF_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R0_INV_0 (.A(tie_lo_T16Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y12__R1_BUF_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R1_INV_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R2_INV_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y12__R2_INV_1 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y12__R3_BUF_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y13__R0_BUF_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R0_INV_0 (.A(tie_lo_T16Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y13__R1_BUF_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R1_INV_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R2_INV_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y13__R2_INV_1 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y13__R3_BUF_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y14__R0_BUF_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R0_INV_0 (.A(tie_lo_T16Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y14__R1_BUF_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R1_INV_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R2_INV_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y14__R2_INV_1 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y14__R3_BUF_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y15__R0_BUF_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R0_INV_0 (.A(tie_lo_T16Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y15__R1_BUF_0 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R1_INV_0 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R2_INV_0 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y15__R2_INV_1 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y15__R3_BUF_0 (.A(tie_lo_T16Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y16__R0_BUF_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R0_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y16__R1_BUF_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R1_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R2_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y16__R2_INV_1 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y16__R3_BUF_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y17__R0_BUF_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R0_INV_0 (.A(tie_lo_T16Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y17__R1_BUF_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R1_INV_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R2_INV_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y17__R2_INV_1 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y17__R3_BUF_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y18__R0_BUF_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R0_INV_0 (.A(tie_lo_T16Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y18__R1_BUF_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R1_INV_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R2_INV_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y18__R2_INV_1 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y18__R3_BUF_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y19__R0_BUF_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R0_INV_0 (.A(tie_lo_T16Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y19__R1_BUF_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R1_INV_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R2_INV_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y19__R2_INV_1 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y19__R3_BUF_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y1__R0_BUF_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R0_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y1__R1_BUF_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R1_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R2_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y1__R2_INV_1 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y1__R3_BUF_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y20__R0_BUF_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R0_INV_0 (.A(tie_lo_T16Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y20__R1_BUF_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R1_INV_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R2_INV_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y20__R2_INV_1 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y20__R3_BUF_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y21__R0_BUF_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R0_INV_0 (.A(tie_lo_T16Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y21__R1_BUF_0 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R1_INV_0 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R2_INV_0 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y21__R2_INV_1 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y21__R3_BUF_0 (.A(tie_lo_T16Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y22__R0_BUF_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R0_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y22__R1_BUF_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R1_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R2_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y22__R2_INV_1 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y22__R3_BUF_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y23__R0_BUF_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R0_INV_0 (.A(tie_lo_T16Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y23__R1_BUF_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R1_INV_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R2_INV_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y23__R2_INV_1 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y23__R3_BUF_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y24__R0_BUF_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R0_INV_0 (.A(tie_lo_T16Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y24__R1_BUF_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R1_INV_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R2_INV_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y24__R2_INV_1 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y24__R3_BUF_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y25__R0_BUF_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R0_INV_0 (.A(tie_lo_T16Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y25__R1_BUF_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R1_INV_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R2_INV_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y25__R2_INV_1 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y25__R3_BUF_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y26__R0_BUF_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R0_INV_0 (.A(tie_lo_T16Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y26__R1_BUF_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R1_INV_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R2_INV_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y26__R2_INV_1 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y26__R3_BUF_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y27__R0_BUF_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R0_INV_0 (.A(tie_lo_T16Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y27__R1_BUF_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R1_INV_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R2_INV_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y27__R2_INV_1 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y27__R3_BUF_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y28__R0_BUF_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R0_INV_0 (.A(tie_lo_T16Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y28__R1_BUF_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R1_INV_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R2_INV_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y28__R2_INV_1 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y28__R3_BUF_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y29__R0_BUF_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R0_INV_0 (.A(tie_lo_T16Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y29__R1_BUF_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R1_INV_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R2_INV_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y29__R2_INV_1 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y29__R3_BUF_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y2__R0_BUF_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R0_INV_0 (.A(tie_lo_T16Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y2__R1_BUF_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R1_INV_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R2_INV_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y2__R2_INV_1 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y2__R3_BUF_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y30__R0_BUF_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R0_INV_0 (.A(tie_lo_T16Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y30__R1_BUF_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R1_INV_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R2_INV_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y30__R2_INV_1 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y30__R3_BUF_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y31__R0_BUF_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R0_INV_0 (.A(tie_lo_T16Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y31__R1_BUF_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R1_INV_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R2_INV_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y31__R2_INV_1 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y31__R3_BUF_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y32__R0_BUF_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R0_INV_0 (.A(tie_lo_T16Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y32__R1_BUF_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R1_INV_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R2_INV_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y32__R2_INV_1 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y32__R3_BUF_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y33__R0_BUF_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R0_INV_0 (.A(tie_lo_T16Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y33__R1_BUF_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R1_INV_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R2_INV_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y33__R2_INV_1 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y33__R3_BUF_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y34__R0_BUF_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R0_INV_0 (.A(tie_lo_T16Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y34__R1_BUF_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R1_INV_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R2_INV_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y34__R2_INV_1 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y34__R3_BUF_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y35__R0_BUF_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R0_INV_0 (.A(tie_lo_T16Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y35__R1_BUF_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R1_INV_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R2_INV_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y35__R2_INV_1 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y35__R3_BUF_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y36__R0_BUF_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R0_INV_0 (.A(tie_lo_T16Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y36__R1_BUF_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R1_INV_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R2_INV_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y36__R2_INV_1 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y36__R3_BUF_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y37__R0_BUF_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R0_INV_0 (.A(tie_lo_T16Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y37__R1_BUF_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R1_INV_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R2_INV_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y37__R2_INV_1 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y37__R3_BUF_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y38__R0_BUF_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R0_INV_0 (.A(tie_lo_T16Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y38__R1_BUF_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R1_INV_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R2_INV_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y38__R2_INV_1 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y38__R3_BUF_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y39__R0_BUF_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R0_INV_0 (.A(tie_lo_T16Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y39__R1_BUF_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R1_INV_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R2_INV_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y39__R2_INV_1 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y39__R3_BUF_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y3__R0_BUF_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R0_INV_0 (.A(tie_lo_T16Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y3__R1_BUF_0 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R1_INV_0 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R2_INV_0 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y3__R2_INV_1 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y3__R3_BUF_0 (.A(tie_lo_T16Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y40__R0_BUF_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R0_INV_0 (.A(tie_lo_T16Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y40__R1_BUF_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R1_INV_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R2_INV_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y40__R2_INV_1 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y40__R3_BUF_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y41__R0_BUF_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R0_INV_0 (.A(tie_lo_T16Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y41__R1_BUF_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R1_INV_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R2_INV_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y41__R2_INV_1 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y41__R3_BUF_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y42__R0_BUF_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R0_INV_0 (.A(tie_lo_T16Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y42__R1_BUF_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R1_INV_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R2_INV_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y42__R2_INV_1 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y42__R3_BUF_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y43__R0_BUF_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R0_INV_0 (.A(tie_lo_T16Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y43__R1_BUF_0 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R1_INV_0 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R2_INV_0 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y43__R2_INV_1 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y43__R3_BUF_0 (.A(tie_lo_T16Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y44__R0_BUF_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R0_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y44__R1_BUF_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R1_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R2_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y44__R2_INV_1 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y44__R3_BUF_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y45__R0_BUF_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R0_INV_0 (.A(tie_lo_T16Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y45__R1_BUF_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R1_INV_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R2_INV_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y45__R2_INV_1 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y45__R3_BUF_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y46__R0_BUF_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R0_INV_0 (.A(tie_lo_T16Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y46__R1_BUF_0 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R1_INV_0 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R2_INV_0 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y46__R2_INV_1 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y46__R3_BUF_0 (.A(tie_lo_T16Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y47__R0_BUF_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R0_INV_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y47__R1_BUF_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R1_INV_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R2_INV_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y47__R2_INV_1 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y47__R3_BUF_0 (.A(tie_lo_T16Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y48__R0_BUF_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R0_INV_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y48__R1_BUF_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R1_INV_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R2_INV_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y48__R2_INV_1 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y48__R3_BUF_0 (.A(tie_lo_T16Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y49__R0_BUF_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R0_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y49__R1_BUF_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R1_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R2_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y49__R2_INV_1 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y49__R3_BUF_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y4__R0_BUF_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R0_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y4__R1_BUF_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R1_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R2_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y4__R2_INV_1 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y4__R3_BUF_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y50__R0_BUF_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R0_INV_0 (.A(tie_lo_T16Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y50__R1_BUF_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R1_INV_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R2_INV_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y50__R2_INV_1 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y50__R3_BUF_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y51__R0_BUF_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R0_INV_0 (.A(tie_lo_T16Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y51__R1_BUF_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R1_INV_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R2_INV_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y51__R2_INV_1 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y51__R3_BUF_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y52__R0_BUF_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R0_INV_0 (.A(tie_lo_T16Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y52__R1_BUF_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R1_INV_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R2_INV_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y52__R2_INV_1 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y52__R3_BUF_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y53__R0_BUF_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R0_INV_0 (.A(tie_lo_T16Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y53__R1_BUF_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R1_INV_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R2_INV_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y53__R2_INV_1 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y53__R3_BUF_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y54__R0_BUF_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R0_INV_0 (.A(tie_lo_T16Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y54__R1_BUF_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R1_INV_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R2_INV_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y54__R2_INV_1 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y54__R3_BUF_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y55__R0_BUF_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R0_INV_0 (.A(tie_lo_T16Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y55__R1_BUF_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R1_INV_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R2_INV_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y55__R2_INV_1 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y55__R3_BUF_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y56__R0_BUF_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R0_INV_0 (.A(tie_lo_T16Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y56__R1_BUF_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R1_INV_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R2_INV_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y56__R2_INV_1 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y56__R3_BUF_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y57__R0_BUF_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R0_INV_0 (.A(tie_lo_T16Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y57__R1_BUF_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R1_INV_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R2_INV_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y57__R2_INV_1 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y57__R3_BUF_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y58__R0_BUF_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R0_INV_0 (.A(tie_lo_T16Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y58__R1_BUF_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R1_INV_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R2_INV_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y58__R2_INV_1 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y58__R3_BUF_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y59__R0_BUF_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R0_INV_0 (.A(tie_lo_T16Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y59__R1_BUF_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R1_INV_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R2_INV_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y59__R2_INV_1 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y59__R3_BUF_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y5__R0_BUF_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R0_INV_0 (.A(tie_lo_T16Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y5__R1_BUF_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R1_INV_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R2_INV_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y5__R2_INV_1 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y5__R3_BUF_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y60__R0_BUF_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R0_INV_0 (.A(tie_lo_T16Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y60__R1_BUF_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R1_INV_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R2_INV_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y60__R2_INV_1 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y60__R3_BUF_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y61__R0_BUF_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R0_INV_0 (.A(tie_lo_T16Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y61__R1_BUF_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R1_INV_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R2_INV_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y61__R2_INV_1 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y61__R3_BUF_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y62__R0_BUF_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R0_INV_0 (.A(tie_lo_T16Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y62__R1_BUF_0 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R1_INV_0 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R2_INV_0 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y62__R2_INV_1 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y62__R3_BUF_0 (.A(tie_lo_T16Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y63__R0_BUF_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R0_INV_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y63__R1_BUF_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R1_INV_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R2_INV_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y63__R2_INV_1 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y63__R3_BUF_0 (.A(tie_lo_T16Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y64__R0_BUF_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R0_INV_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y64__R1_BUF_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R1_INV_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R2_INV_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y64__R2_INV_1 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y64__R3_BUF_0 (.A(tie_lo_T16Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y65__R0_BUF_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R0_INV_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y65__R1_BUF_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R1_INV_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R2_INV_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y65__R2_INV_1 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y65__R3_BUF_0 (.A(tie_lo_T16Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y66__R0_BUF_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R0_INV_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y66__R1_BUF_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R1_INV_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R2_INV_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y66__R2_INV_1 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y66__R3_BUF_0 (.A(tie_lo_T16Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y67__R0_BUF_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R0_INV_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y67__R1_BUF_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R1_INV_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R2_INV_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y67__R2_INV_1 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y67__R3_BUF_0 (.A(tie_lo_T16Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y68__R0_BUF_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R0_INV_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y68__R1_BUF_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R1_INV_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R2_INV_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y68__R2_INV_1 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y68__R3_BUF_0 (.A(tie_lo_T16Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y69__R0_BUF_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R0_INV_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y69__R1_BUF_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R1_INV_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R2_INV_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y69__R2_INV_1 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y69__R3_BUF_0 (.A(tie_lo_T16Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y6__R0_BUF_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R0_INV_0 (.A(tie_lo_T16Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y6__R1_BUF_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R1_INV_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R2_INV_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y6__R2_INV_1 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y6__R3_BUF_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y70__R0_BUF_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R0_INV_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y70__R1_BUF_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R1_INV_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R2_INV_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y70__R2_INV_1 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y70__R3_BUF_0 (.A(tie_lo_T16Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y71__R0_BUF_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R0_INV_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y71__R1_BUF_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R1_INV_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R2_INV_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y71__R2_INV_1 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y71__R3_BUF_0 (.A(tie_lo_T16Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y72__R0_BUF_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R0_INV_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y72__R1_BUF_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R1_INV_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R2_INV_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y72__R2_INV_1 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y72__R3_BUF_0 (.A(tie_lo_T16Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y73__R0_BUF_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R0_INV_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y73__R1_BUF_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R1_INV_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R2_INV_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y73__R2_INV_1 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y73__R3_BUF_0 (.A(tie_lo_T16Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y74__R0_BUF_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R0_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y74__R1_BUF_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R1_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R2_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y74__R2_INV_1 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y74__R3_BUF_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y75__R0_BUF_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R0_INV_0 (.A(tie_lo_T16Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y75__R1_BUF_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R1_INV_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R2_INV_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y75__R2_INV_1 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y75__R3_BUF_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y76__R0_BUF_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R0_INV_0 (.A(tie_lo_T16Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y76__R1_BUF_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R1_INV_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R2_INV_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y76__R2_INV_1 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y76__R3_BUF_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y77__R0_BUF_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R0_INV_0 (.A(tie_lo_T16Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y77__R1_BUF_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R1_INV_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R2_INV_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y77__R2_INV_1 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y77__R3_BUF_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y78__R0_BUF_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R0_INV_0 (.A(tie_lo_T16Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y78__R1_BUF_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R1_INV_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R2_INV_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y78__R2_INV_1 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y78__R3_BUF_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y79__R0_BUF_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R0_INV_0 (.A(tie_lo_T16Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y79__R1_BUF_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R1_INV_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R2_INV_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y79__R2_INV_1 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y79__R3_BUF_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y7__R0_BUF_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R0_INV_0 (.A(tie_lo_T16Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y7__R1_BUF_0 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R1_INV_0 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R2_INV_0 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y7__R2_INV_1 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y7__R3_BUF_0 (.A(tie_lo_T16Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y80__R0_BUF_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R0_INV_0 (.A(tie_lo_T16Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y80__R1_BUF_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R1_INV_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R2_INV_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y80__R2_INV_1 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y80__R3_BUF_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y81__R0_BUF_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R0_INV_0 (.A(tie_lo_T16Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y81__R1_BUF_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R1_INV_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R2_INV_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y81__R2_INV_1 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y81__R3_BUF_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y82__R0_BUF_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R0_INV_0 (.A(tie_lo_T16Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y82__R1_BUF_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R1_INV_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R2_INV_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y82__R2_INV_1 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y82__R3_BUF_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y83__R0_BUF_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R0_INV_0 (.A(tie_lo_T16Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y83__R1_BUF_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R1_INV_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R2_INV_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y83__R2_INV_1 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y83__R3_BUF_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y84__R0_BUF_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R0_INV_0 (.A(tie_lo_T16Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y84__R1_BUF_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R1_INV_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R2_INV_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y84__R2_INV_1 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y84__R3_BUF_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y85__R0_BUF_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R0_INV_0 (.A(tie_lo_T16Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y85__R1_BUF_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R1_INV_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R2_INV_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y85__R2_INV_1 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y85__R3_BUF_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y86__R0_BUF_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R0_INV_0 (.A(tie_lo_T16Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y86__R1_BUF_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R1_INV_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R2_INV_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y86__R2_INV_1 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y86__R3_BUF_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y87__R0_BUF_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R0_INV_0 (.A(tie_lo_T16Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y87__R1_BUF_0 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R1_INV_0 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R2_INV_0 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y87__R2_INV_1 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y87__R3_BUF_0 (.A(tie_lo_T16Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y88__R0_BUF_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R0_INV_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y88__R1_BUF_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R1_INV_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R2_INV_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y88__R2_INV_1 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y88__R3_BUF_0 (.A(tie_lo_T16Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y89__R0_BUF_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R0_INV_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y89__R1_BUF_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R1_INV_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R2_INV_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y89__R2_INV_1 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y89__R3_BUF_0 (.A(tie_lo_T16Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y8__R0_BUF_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R0_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y8__R1_BUF_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R1_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R2_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y8__R2_INV_1 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y8__R3_BUF_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y9__R0_BUF_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R0_INV_0 (.A(tie_lo_T16Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y9__R1_BUF_0 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R1_INV_0 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T16Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R2_INV_0 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T16Y9__R2_INV_1 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T16Y9__R3_BUF_0 (.A(tie_lo_T16Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y0__R0_BUF_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R0_INV_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y0__R1_BUF_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R1_INV_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R2_INV_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y0__R2_INV_1 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y0__R3_BUF_0 (.A(tie_lo_T17Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y10__R0_BUF_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R0_INV_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y10__R1_BUF_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R1_INV_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R2_INV_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y10__R2_INV_1 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y10__R3_BUF_0 (.A(tie_lo_T17Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y11__R0_BUF_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R0_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y11__R1_BUF_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R1_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R2_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y11__R2_INV_1 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y11__R3_BUF_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y12__R0_BUF_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R0_INV_0 (.A(tie_lo_T17Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y12__R1_BUF_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R1_INV_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R2_INV_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y12__R2_INV_1 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y12__R3_BUF_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y13__R0_BUF_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R0_INV_0 (.A(tie_lo_T17Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y13__R1_BUF_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R1_INV_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R2_INV_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y13__R2_INV_1 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y13__R3_BUF_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y14__R0_BUF_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R0_INV_0 (.A(tie_lo_T17Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y14__R1_BUF_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R1_INV_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R2_INV_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y14__R2_INV_1 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y14__R3_BUF_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y15__R0_BUF_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R0_INV_0 (.A(tie_lo_T17Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y15__R1_BUF_0 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R1_INV_0 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R2_INV_0 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y15__R2_INV_1 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y15__R3_BUF_0 (.A(tie_lo_T17Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y16__R0_BUF_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R0_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y16__R1_BUF_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R1_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R2_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y16__R2_INV_1 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y16__R3_BUF_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y17__R0_BUF_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R0_INV_0 (.A(tie_lo_T17Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y17__R1_BUF_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R1_INV_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R2_INV_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y17__R2_INV_1 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y17__R3_BUF_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y18__R0_BUF_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R0_INV_0 (.A(tie_lo_T17Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y18__R1_BUF_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R1_INV_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R2_INV_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y18__R2_INV_1 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y18__R3_BUF_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y19__R0_BUF_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R0_INV_0 (.A(tie_lo_T17Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y19__R1_BUF_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R1_INV_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R2_INV_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y19__R2_INV_1 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y19__R3_BUF_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y1__R0_BUF_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R0_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y1__R1_BUF_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R1_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R2_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y1__R2_INV_1 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y1__R3_BUF_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y20__R0_BUF_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R0_INV_0 (.A(tie_lo_T17Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y20__R1_BUF_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R1_INV_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R2_INV_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y20__R2_INV_1 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y20__R3_BUF_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y21__R0_BUF_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R0_INV_0 (.A(tie_lo_T17Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y21__R1_BUF_0 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R1_INV_0 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R2_INV_0 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y21__R2_INV_1 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y21__R3_BUF_0 (.A(tie_lo_T17Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y22__R0_BUF_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R0_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y22__R1_BUF_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R1_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R2_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y22__R2_INV_1 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y22__R3_BUF_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y23__R0_BUF_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R0_INV_0 (.A(tie_lo_T17Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y23__R1_BUF_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R1_INV_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R2_INV_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y23__R2_INV_1 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y23__R3_BUF_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y24__R0_BUF_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R0_INV_0 (.A(tie_lo_T17Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y24__R1_BUF_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R1_INV_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R2_INV_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y24__R2_INV_1 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y24__R3_BUF_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y25__R0_BUF_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R0_INV_0 (.A(tie_lo_T17Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y25__R1_BUF_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R1_INV_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R2_INV_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y25__R2_INV_1 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y25__R3_BUF_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y26__R0_BUF_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R0_INV_0 (.A(tie_lo_T17Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y26__R1_BUF_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R1_INV_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R2_INV_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y26__R2_INV_1 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y26__R3_BUF_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y27__R0_BUF_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R0_INV_0 (.A(tie_lo_T17Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y27__R1_BUF_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R1_INV_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R2_INV_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y27__R2_INV_1 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y27__R3_BUF_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y28__R0_BUF_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R0_INV_0 (.A(tie_lo_T17Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y28__R1_BUF_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R1_INV_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R2_INV_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y28__R2_INV_1 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y28__R3_BUF_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y29__R0_BUF_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R0_INV_0 (.A(tie_lo_T17Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y29__R1_BUF_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R1_INV_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R2_INV_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y29__R2_INV_1 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y29__R3_BUF_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y2__R0_BUF_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R0_INV_0 (.A(tie_lo_T17Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y2__R1_BUF_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R1_INV_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R2_INV_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y2__R2_INV_1 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y2__R3_BUF_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y30__R0_BUF_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R0_INV_0 (.A(tie_lo_T17Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y30__R1_BUF_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R1_INV_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R2_INV_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y30__R2_INV_1 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y30__R3_BUF_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y31__R0_BUF_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R0_INV_0 (.A(tie_lo_T17Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y31__R1_BUF_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R1_INV_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R2_INV_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y31__R2_INV_1 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y31__R3_BUF_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y32__R0_BUF_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R0_INV_0 (.A(tie_lo_T17Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y32__R1_BUF_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R1_INV_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R2_INV_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y32__R2_INV_1 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y32__R3_BUF_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y33__R0_BUF_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R0_INV_0 (.A(tie_lo_T17Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y33__R1_BUF_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R1_INV_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R2_INV_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y33__R2_INV_1 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y33__R3_BUF_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y34__R0_BUF_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R0_INV_0 (.A(tie_lo_T17Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y34__R1_BUF_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R1_INV_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R2_INV_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y34__R2_INV_1 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y34__R3_BUF_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y35__R0_BUF_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R0_INV_0 (.A(tie_lo_T17Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y35__R1_BUF_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R1_INV_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R2_INV_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y35__R2_INV_1 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y35__R3_BUF_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y36__R0_BUF_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R0_INV_0 (.A(tie_lo_T17Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y36__R1_BUF_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R1_INV_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R2_INV_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y36__R2_INV_1 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y36__R3_BUF_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y37__R0_BUF_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R0_INV_0 (.A(tie_lo_T17Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y37__R1_BUF_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R1_INV_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R2_INV_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y37__R2_INV_1 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y37__R3_BUF_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y38__R0_BUF_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R0_INV_0 (.A(tie_lo_T17Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y38__R1_BUF_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R1_INV_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R2_INV_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y38__R2_INV_1 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y38__R3_BUF_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y39__R0_BUF_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R0_INV_0 (.A(tie_lo_T17Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y39__R1_BUF_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R1_INV_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R2_INV_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y39__R2_INV_1 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y39__R3_BUF_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y3__R0_BUF_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R0_INV_0 (.A(tie_lo_T17Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y3__R1_BUF_0 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R1_INV_0 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R2_INV_0 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y3__R2_INV_1 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y3__R3_BUF_0 (.A(tie_lo_T17Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y40__R0_BUF_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R0_INV_0 (.A(tie_lo_T17Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y40__R1_BUF_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R1_INV_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R2_INV_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y40__R2_INV_1 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y40__R3_BUF_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y41__R0_BUF_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R0_INV_0 (.A(tie_lo_T17Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y41__R1_BUF_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R1_INV_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R2_INV_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y41__R2_INV_1 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y41__R3_BUF_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y42__R0_BUF_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R0_INV_0 (.A(tie_lo_T17Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y42__R1_BUF_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R1_INV_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R2_INV_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y42__R2_INV_1 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y42__R3_BUF_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y43__R0_BUF_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R0_INV_0 (.A(tie_lo_T17Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y43__R1_BUF_0 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R1_INV_0 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R2_INV_0 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y43__R2_INV_1 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y43__R3_BUF_0 (.A(tie_lo_T17Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y44__R0_BUF_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R0_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y44__R1_BUF_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R1_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R2_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y44__R2_INV_1 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y44__R3_BUF_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y45__R0_BUF_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R0_INV_0 (.A(tie_lo_T17Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y45__R1_BUF_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R1_INV_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R2_INV_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y45__R2_INV_1 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y45__R3_BUF_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y46__R0_BUF_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R0_INV_0 (.A(tie_lo_T17Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y46__R1_BUF_0 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R1_INV_0 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R2_INV_0 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y46__R2_INV_1 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y46__R3_BUF_0 (.A(tie_lo_T17Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y47__R0_BUF_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R0_INV_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y47__R1_BUF_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R1_INV_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R2_INV_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y47__R2_INV_1 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y47__R3_BUF_0 (.A(tie_lo_T17Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y48__R0_BUF_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R0_INV_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y48__R1_BUF_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R1_INV_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R2_INV_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y48__R2_INV_1 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y48__R3_BUF_0 (.A(tie_lo_T17Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y49__R0_BUF_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R0_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y49__R1_BUF_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R1_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R2_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y49__R2_INV_1 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y49__R3_BUF_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y4__R0_BUF_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R0_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y4__R1_BUF_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R1_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R2_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y4__R2_INV_1 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y4__R3_BUF_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y50__R0_BUF_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R0_INV_0 (.A(tie_lo_T17Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y50__R1_BUF_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R1_INV_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R2_INV_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y50__R2_INV_1 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y50__R3_BUF_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y51__R0_BUF_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R0_INV_0 (.A(tie_lo_T17Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y51__R1_BUF_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R1_INV_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R2_INV_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y51__R2_INV_1 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y51__R3_BUF_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y52__R0_BUF_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R0_INV_0 (.A(tie_lo_T17Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y52__R1_BUF_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R1_INV_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R2_INV_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y52__R2_INV_1 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y52__R3_BUF_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y53__R0_BUF_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R0_INV_0 (.A(tie_lo_T17Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y53__R1_BUF_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R1_INV_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R2_INV_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y53__R2_INV_1 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y53__R3_BUF_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y54__R0_BUF_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R0_INV_0 (.A(tie_lo_T17Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y54__R1_BUF_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R1_INV_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R2_INV_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y54__R2_INV_1 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y54__R3_BUF_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y55__R0_BUF_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R0_INV_0 (.A(tie_lo_T17Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y55__R1_BUF_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R1_INV_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R2_INV_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y55__R2_INV_1 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y55__R3_BUF_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y56__R0_BUF_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R0_INV_0 (.A(tie_lo_T17Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y56__R1_BUF_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R1_INV_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R2_INV_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y56__R2_INV_1 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y56__R3_BUF_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y57__R0_BUF_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R0_INV_0 (.A(tie_lo_T17Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y57__R1_BUF_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R1_INV_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R2_INV_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y57__R2_INV_1 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y57__R3_BUF_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y58__R0_BUF_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R0_INV_0 (.A(tie_lo_T17Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y58__R1_BUF_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R1_INV_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R2_INV_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y58__R2_INV_1 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y58__R3_BUF_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y59__R0_BUF_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R0_INV_0 (.A(tie_lo_T17Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y59__R1_BUF_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R1_INV_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R2_INV_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y59__R2_INV_1 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y59__R3_BUF_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y5__R0_BUF_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R0_INV_0 (.A(tie_lo_T17Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y5__R1_BUF_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R1_INV_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R2_INV_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y5__R2_INV_1 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y5__R3_BUF_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y60__R0_BUF_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R0_INV_0 (.A(tie_lo_T17Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y60__R1_BUF_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R1_INV_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R2_INV_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y60__R2_INV_1 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y60__R3_BUF_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y61__R0_BUF_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R0_INV_0 (.A(tie_lo_T17Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y61__R1_BUF_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R1_INV_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R2_INV_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y61__R2_INV_1 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y61__R3_BUF_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y62__R0_BUF_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R0_INV_0 (.A(tie_lo_T17Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y62__R1_BUF_0 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R1_INV_0 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R2_INV_0 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y62__R2_INV_1 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y62__R3_BUF_0 (.A(tie_lo_T17Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y63__R0_BUF_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R0_INV_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y63__R1_BUF_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R1_INV_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R2_INV_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y63__R2_INV_1 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y63__R3_BUF_0 (.A(tie_lo_T17Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y64__R0_BUF_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R0_INV_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y64__R1_BUF_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R1_INV_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R2_INV_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y64__R2_INV_1 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y64__R3_BUF_0 (.A(tie_lo_T17Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y65__R0_BUF_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R0_INV_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y65__R1_BUF_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R1_INV_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R2_INV_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y65__R2_INV_1 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y65__R3_BUF_0 (.A(tie_lo_T17Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y66__R0_BUF_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R0_INV_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y66__R1_BUF_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R1_INV_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R2_INV_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y66__R2_INV_1 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y66__R3_BUF_0 (.A(tie_lo_T17Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y67__R0_BUF_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R0_INV_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y67__R1_BUF_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R1_INV_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R2_INV_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y67__R2_INV_1 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y67__R3_BUF_0 (.A(tie_lo_T17Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y68__R0_BUF_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R0_INV_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y68__R1_BUF_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R1_INV_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R2_INV_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y68__R2_INV_1 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y68__R3_BUF_0 (.A(tie_lo_T17Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y69__R0_BUF_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R0_INV_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y69__R1_BUF_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R1_INV_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R2_INV_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y69__R2_INV_1 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y69__R3_BUF_0 (.A(tie_lo_T17Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y6__R0_BUF_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R0_INV_0 (.A(tie_lo_T17Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y6__R1_BUF_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R1_INV_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R2_INV_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y6__R2_INV_1 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y6__R3_BUF_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y70__R0_BUF_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R0_INV_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y70__R1_BUF_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R1_INV_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R2_INV_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y70__R2_INV_1 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y70__R3_BUF_0 (.A(tie_lo_T17Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y71__R0_BUF_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R0_INV_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y71__R1_BUF_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R1_INV_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R2_INV_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y71__R2_INV_1 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y71__R3_BUF_0 (.A(tie_lo_T17Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y72__R0_BUF_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R0_INV_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y72__R1_BUF_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R1_INV_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R2_INV_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y72__R2_INV_1 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y72__R3_BUF_0 (.A(tie_lo_T17Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y73__R0_BUF_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R0_INV_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y73__R1_BUF_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R1_INV_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R2_INV_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y73__R2_INV_1 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y73__R3_BUF_0 (.A(tie_lo_T17Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y74__R0_BUF_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R0_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y74__R1_BUF_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R1_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R2_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y74__R2_INV_1 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y74__R3_BUF_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y75__R0_BUF_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R0_INV_0 (.A(tie_lo_T17Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y75__R1_BUF_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R1_INV_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R2_INV_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y75__R2_INV_1 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y75__R3_BUF_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y76__R0_BUF_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R0_INV_0 (.A(tie_lo_T17Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y76__R1_BUF_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R1_INV_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R2_INV_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y76__R2_INV_1 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y76__R3_BUF_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y77__R0_BUF_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R0_INV_0 (.A(tie_lo_T17Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y77__R1_BUF_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R1_INV_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R2_INV_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y77__R2_INV_1 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y77__R3_BUF_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y78__R0_BUF_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R0_INV_0 (.A(tie_lo_T17Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y78__R1_BUF_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R1_INV_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R2_INV_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y78__R2_INV_1 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y78__R3_BUF_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y79__R0_BUF_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R0_INV_0 (.A(tie_lo_T17Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y79__R1_BUF_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R1_INV_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R2_INV_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y79__R2_INV_1 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y79__R3_BUF_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y7__R0_BUF_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R0_INV_0 (.A(tie_lo_T17Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y7__R1_BUF_0 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R1_INV_0 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R2_INV_0 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y7__R2_INV_1 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y7__R3_BUF_0 (.A(tie_lo_T17Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y80__R0_BUF_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R0_INV_0 (.A(tie_lo_T17Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y80__R1_BUF_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R1_INV_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R2_INV_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y80__R2_INV_1 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y80__R3_BUF_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y81__R0_BUF_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R0_INV_0 (.A(tie_lo_T17Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y81__R1_BUF_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R1_INV_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R2_INV_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y81__R2_INV_1 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y81__R3_BUF_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y82__R0_BUF_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R0_INV_0 (.A(tie_lo_T17Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y82__R1_BUF_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R1_INV_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R2_INV_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y82__R2_INV_1 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y82__R3_BUF_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y83__R0_BUF_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R0_INV_0 (.A(tie_lo_T17Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y83__R1_BUF_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R1_INV_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R2_INV_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y83__R2_INV_1 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y83__R3_BUF_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y84__R0_BUF_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R0_INV_0 (.A(tie_lo_T17Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y84__R1_BUF_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R1_INV_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R2_INV_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y84__R2_INV_1 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y84__R3_BUF_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y85__R0_BUF_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R0_INV_0 (.A(tie_lo_T17Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y85__R1_BUF_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R1_INV_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R2_INV_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y85__R2_INV_1 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y85__R3_BUF_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y86__R0_BUF_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R0_INV_0 (.A(tie_lo_T17Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y86__R1_BUF_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R1_INV_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R2_INV_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y86__R2_INV_1 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y86__R3_BUF_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y87__R0_BUF_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R0_INV_0 (.A(tie_lo_T17Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y87__R1_BUF_0 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R1_INV_0 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R2_INV_0 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y87__R2_INV_1 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y87__R3_BUF_0 (.A(tie_lo_T17Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y88__R0_BUF_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R0_INV_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y88__R1_BUF_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R1_INV_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R2_INV_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y88__R2_INV_1 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y88__R3_BUF_0 (.A(tie_lo_T17Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y89__R0_BUF_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R0_INV_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y89__R1_BUF_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R1_INV_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R2_INV_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y89__R2_INV_1 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y89__R3_BUF_0 (.A(tie_lo_T17Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y8__R0_BUF_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R0_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y8__R1_BUF_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R1_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R2_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y8__R2_INV_1 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y8__R3_BUF_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y9__R0_BUF_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R0_INV_0 (.A(tie_lo_T17Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y9__R1_BUF_0 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R1_INV_0 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T17Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R2_INV_0 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T17Y9__R2_INV_1 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T17Y9__R3_BUF_0 (.A(tie_lo_T17Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y0__R0_BUF_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R0_INV_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y0__R1_BUF_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R1_INV_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R2_INV_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y0__R2_INV_1 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y0__R3_BUF_0 (.A(tie_lo_T18Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y10__R0_BUF_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R0_INV_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y10__R1_BUF_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R1_INV_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R2_INV_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y10__R2_INV_1 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y10__R3_BUF_0 (.A(tie_lo_T18Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y11__R0_BUF_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R0_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y11__R1_BUF_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R1_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R2_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y11__R2_INV_1 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y11__R3_BUF_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y12__R0_BUF_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R0_INV_0 (.A(tie_lo_T18Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y12__R1_BUF_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R1_INV_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R2_INV_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y12__R2_INV_1 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y12__R3_BUF_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y13__R0_BUF_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R0_INV_0 (.A(tie_lo_T18Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y13__R1_BUF_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R1_INV_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R2_INV_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y13__R2_INV_1 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y13__R3_BUF_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y14__R0_BUF_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R0_INV_0 (.A(tie_lo_T18Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y14__R1_BUF_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R1_INV_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R2_INV_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y14__R2_INV_1 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y14__R3_BUF_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y15__R0_BUF_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R0_INV_0 (.A(tie_lo_T18Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y15__R1_BUF_0 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R1_INV_0 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R2_INV_0 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y15__R2_INV_1 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y15__R3_BUF_0 (.A(tie_lo_T18Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y16__R0_BUF_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R0_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y16__R1_BUF_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R1_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R2_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y16__R2_INV_1 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y16__R3_BUF_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y17__R0_BUF_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R0_INV_0 (.A(tie_lo_T18Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y17__R1_BUF_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R1_INV_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R2_INV_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y17__R2_INV_1 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y17__R3_BUF_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y18__R0_BUF_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R0_INV_0 (.A(tie_lo_T18Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y18__R1_BUF_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R1_INV_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R2_INV_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y18__R2_INV_1 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y18__R3_BUF_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y19__R0_BUF_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R0_INV_0 (.A(tie_lo_T18Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y19__R1_BUF_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R1_INV_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R2_INV_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y19__R2_INV_1 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y19__R3_BUF_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y1__R0_BUF_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R0_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y1__R1_BUF_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R1_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R2_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y1__R2_INV_1 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y1__R3_BUF_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y20__R0_BUF_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R0_INV_0 (.A(tie_lo_T18Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y20__R1_BUF_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R1_INV_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R2_INV_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y20__R2_INV_1 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y20__R3_BUF_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y21__R0_BUF_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R0_INV_0 (.A(tie_lo_T18Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y21__R1_BUF_0 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R1_INV_0 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R2_INV_0 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y21__R2_INV_1 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y21__R3_BUF_0 (.A(tie_lo_T18Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y22__R0_BUF_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R0_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y22__R1_BUF_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R1_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R2_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y22__R2_INV_1 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y22__R3_BUF_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y23__R0_BUF_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R0_INV_0 (.A(tie_lo_T18Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y23__R1_BUF_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R1_INV_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R2_INV_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y23__R2_INV_1 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y23__R3_BUF_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y24__R0_BUF_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R0_INV_0 (.A(tie_lo_T18Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y24__R1_BUF_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R1_INV_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R2_INV_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y24__R2_INV_1 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y24__R3_BUF_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y25__R0_BUF_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R0_INV_0 (.A(tie_lo_T18Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y25__R1_BUF_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R1_INV_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R2_INV_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y25__R2_INV_1 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y25__R3_BUF_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y26__R0_BUF_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R0_INV_0 (.A(tie_lo_T18Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y26__R1_BUF_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R1_INV_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R2_INV_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y26__R2_INV_1 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y26__R3_BUF_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y27__R0_BUF_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R0_INV_0 (.A(tie_lo_T18Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y27__R1_BUF_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R1_INV_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R2_INV_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y27__R2_INV_1 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y27__R3_BUF_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y28__R0_BUF_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R0_INV_0 (.A(tie_lo_T18Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y28__R1_BUF_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R1_INV_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R2_INV_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y28__R2_INV_1 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y28__R3_BUF_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y29__R0_BUF_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R0_INV_0 (.A(tie_lo_T18Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y29__R1_BUF_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R1_INV_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R2_INV_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y29__R2_INV_1 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y29__R3_BUF_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y2__R0_BUF_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R0_INV_0 (.A(tie_lo_T18Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y2__R1_BUF_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R1_INV_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R2_INV_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y2__R2_INV_1 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y2__R3_BUF_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y30__R0_BUF_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R0_INV_0 (.A(tie_lo_T18Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y30__R1_BUF_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R1_INV_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R2_INV_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y30__R2_INV_1 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y30__R3_BUF_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y31__R0_BUF_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R0_INV_0 (.A(tie_lo_T18Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y31__R1_BUF_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R1_INV_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R2_INV_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y31__R2_INV_1 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y31__R3_BUF_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y32__R0_BUF_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R0_INV_0 (.A(tie_lo_T18Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y32__R1_BUF_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R1_INV_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R2_INV_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y32__R2_INV_1 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y32__R3_BUF_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y33__R0_BUF_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R0_INV_0 (.A(tie_lo_T18Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y33__R1_BUF_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R1_INV_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R2_INV_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y33__R2_INV_1 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y33__R3_BUF_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y34__R0_BUF_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R0_INV_0 (.A(tie_lo_T18Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y34__R1_BUF_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R1_INV_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R2_INV_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y34__R2_INV_1 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y34__R3_BUF_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y35__R0_BUF_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R0_INV_0 (.A(tie_lo_T18Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y35__R1_BUF_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R1_INV_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R2_INV_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y35__R2_INV_1 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y35__R3_BUF_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y36__R0_BUF_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R0_INV_0 (.A(tie_lo_T18Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y36__R1_BUF_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R1_INV_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R2_INV_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y36__R2_INV_1 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y36__R3_BUF_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y37__R0_BUF_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R0_INV_0 (.A(tie_lo_T18Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y37__R1_BUF_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R1_INV_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R2_INV_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y37__R2_INV_1 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y37__R3_BUF_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y38__R0_BUF_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R0_INV_0 (.A(tie_lo_T18Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y38__R1_BUF_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R1_INV_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R2_INV_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y38__R2_INV_1 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y38__R3_BUF_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y39__R0_BUF_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R0_INV_0 (.A(tie_lo_T18Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y39__R1_BUF_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R1_INV_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R2_INV_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y39__R2_INV_1 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y39__R3_BUF_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y3__R0_BUF_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R0_INV_0 (.A(tie_lo_T18Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y3__R1_BUF_0 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R1_INV_0 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R2_INV_0 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y3__R2_INV_1 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y3__R3_BUF_0 (.A(tie_lo_T18Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y40__R0_BUF_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R0_INV_0 (.A(tie_lo_T18Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y40__R1_BUF_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R1_INV_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R2_INV_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y40__R2_INV_1 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y40__R3_BUF_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y41__R0_BUF_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R0_INV_0 (.A(tie_lo_T18Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y41__R1_BUF_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R1_INV_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R2_INV_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y41__R2_INV_1 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y41__R3_BUF_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y42__R0_BUF_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R0_INV_0 (.A(tie_lo_T18Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y42__R1_BUF_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R1_INV_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R2_INV_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y42__R2_INV_1 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y42__R3_BUF_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y43__R0_BUF_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R0_INV_0 (.A(tie_lo_T18Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y43__R1_BUF_0 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R1_INV_0 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R2_INV_0 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y43__R2_INV_1 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y43__R3_BUF_0 (.A(tie_lo_T18Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y44__R0_BUF_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R0_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y44__R1_BUF_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R1_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R2_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y44__R2_INV_1 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y44__R3_BUF_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y45__R0_BUF_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R0_INV_0 (.A(tie_lo_T18Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y45__R1_BUF_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R1_INV_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R2_INV_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y45__R2_INV_1 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y45__R3_BUF_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y46__R0_BUF_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R0_INV_0 (.A(tie_lo_T18Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y46__R1_BUF_0 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R1_INV_0 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R2_INV_0 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y46__R2_INV_1 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y46__R3_BUF_0 (.A(tie_lo_T18Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y47__R0_BUF_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R0_INV_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y47__R1_BUF_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R1_INV_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R2_INV_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y47__R2_INV_1 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y47__R3_BUF_0 (.A(tie_lo_T18Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y48__R0_BUF_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R0_INV_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y48__R1_BUF_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R1_INV_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R2_INV_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y48__R2_INV_1 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y48__R3_BUF_0 (.A(tie_lo_T18Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y49__R0_BUF_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R0_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y49__R1_BUF_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R1_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R2_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y49__R2_INV_1 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y49__R3_BUF_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y4__R0_BUF_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R0_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y4__R1_BUF_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R1_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R2_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y4__R2_INV_1 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y4__R3_BUF_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y50__R0_BUF_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R0_INV_0 (.A(tie_lo_T18Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y50__R1_BUF_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R1_INV_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R2_INV_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y50__R2_INV_1 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y50__R3_BUF_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y51__R0_BUF_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R0_INV_0 (.A(tie_lo_T18Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y51__R1_BUF_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R1_INV_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R2_INV_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y51__R2_INV_1 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y51__R3_BUF_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y52__R0_BUF_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R0_INV_0 (.A(tie_lo_T18Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y52__R1_BUF_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R1_INV_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R2_INV_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y52__R2_INV_1 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y52__R3_BUF_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y53__R0_BUF_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R0_INV_0 (.A(tie_lo_T18Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y53__R1_BUF_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R1_INV_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R2_INV_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y53__R2_INV_1 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y53__R3_BUF_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y54__R0_BUF_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R0_INV_0 (.A(tie_lo_T18Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y54__R1_BUF_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R1_INV_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R2_INV_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y54__R2_INV_1 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y54__R3_BUF_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y55__R0_BUF_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R0_INV_0 (.A(tie_lo_T18Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y55__R1_BUF_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R1_INV_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R2_INV_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y55__R2_INV_1 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y55__R3_BUF_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y56__R0_BUF_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R0_INV_0 (.A(tie_lo_T18Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y56__R1_BUF_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R1_INV_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R2_INV_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y56__R2_INV_1 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y56__R3_BUF_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y57__R0_BUF_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R0_INV_0 (.A(tie_lo_T18Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y57__R1_BUF_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R1_INV_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R2_INV_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y57__R2_INV_1 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y57__R3_BUF_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y58__R0_BUF_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R0_INV_0 (.A(tie_lo_T18Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y58__R1_BUF_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R1_INV_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R2_INV_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y58__R2_INV_1 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y58__R3_BUF_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y59__R0_BUF_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R0_INV_0 (.A(tie_lo_T18Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y59__R1_BUF_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R1_INV_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R2_INV_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y59__R2_INV_1 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y59__R3_BUF_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y5__R0_BUF_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R0_INV_0 (.A(tie_lo_T18Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y5__R1_BUF_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R1_INV_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R2_INV_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y5__R2_INV_1 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y5__R3_BUF_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y60__R0_BUF_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R0_INV_0 (.A(tie_lo_T18Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y60__R1_BUF_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R1_INV_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R2_INV_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y60__R2_INV_1 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y60__R3_BUF_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y61__R0_BUF_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R0_INV_0 (.A(tie_lo_T18Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y61__R1_BUF_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R1_INV_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R2_INV_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y61__R2_INV_1 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y61__R3_BUF_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y62__R0_BUF_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R0_INV_0 (.A(tie_lo_T18Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y62__R1_BUF_0 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R1_INV_0 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R2_INV_0 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y62__R2_INV_1 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y62__R3_BUF_0 (.A(tie_lo_T18Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y63__R0_BUF_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R0_INV_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y63__R1_BUF_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R1_INV_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R2_INV_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y63__R2_INV_1 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y63__R3_BUF_0 (.A(tie_lo_T18Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y64__R0_BUF_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R0_INV_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y64__R1_BUF_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R1_INV_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R2_INV_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y64__R2_INV_1 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y64__R3_BUF_0 (.A(tie_lo_T18Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y65__R0_BUF_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R0_INV_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y65__R1_BUF_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R1_INV_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R2_INV_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y65__R2_INV_1 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y65__R3_BUF_0 (.A(tie_lo_T18Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y66__R0_BUF_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R0_INV_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y66__R1_BUF_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R1_INV_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R2_INV_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y66__R2_INV_1 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y66__R3_BUF_0 (.A(tie_lo_T18Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y67__R0_BUF_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R0_INV_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y67__R1_BUF_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R1_INV_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R2_INV_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y67__R2_INV_1 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y67__R3_BUF_0 (.A(tie_lo_T18Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y68__R0_BUF_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R0_INV_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y68__R1_BUF_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R1_INV_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R2_INV_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y68__R2_INV_1 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y68__R3_BUF_0 (.A(tie_lo_T18Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y69__R0_BUF_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R0_INV_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y69__R1_BUF_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R1_INV_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R2_INV_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y69__R2_INV_1 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y69__R3_BUF_0 (.A(tie_lo_T18Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y6__R0_BUF_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R0_INV_0 (.A(tie_lo_T18Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y6__R1_BUF_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R1_INV_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R2_INV_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y6__R2_INV_1 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y6__R3_BUF_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y70__R0_BUF_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R0_INV_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y70__R1_BUF_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R1_INV_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R2_INV_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y70__R2_INV_1 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y70__R3_BUF_0 (.A(tie_lo_T18Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y71__R0_BUF_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R0_INV_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y71__R1_BUF_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R1_INV_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R2_INV_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y71__R2_INV_1 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y71__R3_BUF_0 (.A(tie_lo_T18Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y72__R0_BUF_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R0_INV_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y72__R1_BUF_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R1_INV_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R2_INV_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y72__R2_INV_1 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y72__R3_BUF_0 (.A(tie_lo_T18Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y73__R0_BUF_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R0_INV_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y73__R1_BUF_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R1_INV_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R2_INV_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y73__R2_INV_1 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y73__R3_BUF_0 (.A(tie_lo_T18Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y74__R0_BUF_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R0_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y74__R1_BUF_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R1_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R2_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y74__R2_INV_1 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y74__R3_BUF_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y75__R0_BUF_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R0_INV_0 (.A(tie_lo_T18Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y75__R1_BUF_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R1_INV_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R2_INV_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y75__R2_INV_1 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y75__R3_BUF_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y76__R0_BUF_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R0_INV_0 (.A(tie_lo_T18Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y76__R1_BUF_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R1_INV_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R2_INV_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y76__R2_INV_1 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y76__R3_BUF_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y77__R0_BUF_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R0_INV_0 (.A(tie_lo_T18Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y77__R1_BUF_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R1_INV_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R2_INV_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y77__R2_INV_1 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y77__R3_BUF_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y78__R0_BUF_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R0_INV_0 (.A(tie_lo_T18Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y78__R1_BUF_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R1_INV_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R2_INV_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y78__R2_INV_1 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y78__R3_BUF_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y79__R0_BUF_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R0_INV_0 (.A(tie_lo_T18Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y79__R1_BUF_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R1_INV_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R2_INV_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y79__R2_INV_1 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y79__R3_BUF_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y7__R0_BUF_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R0_INV_0 (.A(tie_lo_T18Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y7__R1_BUF_0 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R1_INV_0 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R2_INV_0 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y7__R2_INV_1 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y7__R3_BUF_0 (.A(tie_lo_T18Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y80__R0_BUF_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R0_INV_0 (.A(tie_lo_T18Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y80__R1_BUF_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R1_INV_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R2_INV_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y80__R2_INV_1 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y80__R3_BUF_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y81__R0_BUF_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R0_INV_0 (.A(tie_lo_T18Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y81__R1_BUF_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R1_INV_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R2_INV_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y81__R2_INV_1 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y81__R3_BUF_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y82__R0_BUF_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R0_INV_0 (.A(tie_lo_T18Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y82__R1_BUF_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R1_INV_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R2_INV_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y82__R2_INV_1 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y82__R3_BUF_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y83__R0_BUF_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R0_INV_0 (.A(tie_lo_T18Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y83__R1_BUF_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R1_INV_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R2_INV_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y83__R2_INV_1 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y83__R3_BUF_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y84__R0_BUF_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R0_INV_0 (.A(tie_lo_T18Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y84__R1_BUF_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R1_INV_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R2_INV_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y84__R2_INV_1 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y84__R3_BUF_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y85__R0_BUF_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R0_INV_0 (.A(tie_lo_T18Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y85__R1_BUF_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R1_INV_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R2_INV_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y85__R2_INV_1 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y85__R3_BUF_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y86__R0_BUF_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R0_INV_0 (.A(tie_lo_T18Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y86__R1_BUF_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R1_INV_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R2_INV_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y86__R2_INV_1 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y86__R3_BUF_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y87__R0_BUF_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R0_INV_0 (.A(tie_lo_T18Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y87__R1_BUF_0 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R1_INV_0 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R2_INV_0 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y87__R2_INV_1 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y87__R3_BUF_0 (.A(tie_lo_T18Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y88__R0_BUF_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R0_INV_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y88__R1_BUF_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R1_INV_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R2_INV_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y88__R2_INV_1 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y88__R3_BUF_0 (.A(tie_lo_T18Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y89__R0_BUF_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R0_INV_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y89__R1_BUF_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R1_INV_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R2_INV_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y89__R2_INV_1 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y89__R3_BUF_0 (.A(tie_lo_T18Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y8__R0_BUF_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R0_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y8__R1_BUF_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R1_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R2_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y8__R2_INV_1 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y8__R3_BUF_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y9__R0_BUF_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R0_INV_0 (.A(tie_lo_T18Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y9__R1_BUF_0 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R1_INV_0 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T18Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R2_INV_0 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T18Y9__R2_INV_1 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T18Y9__R3_BUF_0 (.A(tie_lo_T18Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y0__R0_BUF_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R0_INV_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y0__R1_BUF_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R1_INV_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R2_INV_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y0__R2_INV_1 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y0__R3_BUF_0 (.A(tie_lo_T19Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y10__R0_BUF_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R0_INV_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y10__R1_BUF_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R1_INV_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R2_INV_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y10__R2_INV_1 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y10__R3_BUF_0 (.A(tie_lo_T19Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y11__R0_BUF_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R0_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y11__R1_BUF_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R1_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R2_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y11__R2_INV_1 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y11__R3_BUF_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y12__R0_BUF_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R0_INV_0 (.A(tie_lo_T19Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y12__R1_BUF_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R1_INV_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R2_INV_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y12__R2_INV_1 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y12__R3_BUF_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y13__R0_BUF_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R0_INV_0 (.A(tie_lo_T19Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y13__R1_BUF_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R1_INV_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R2_INV_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y13__R2_INV_1 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y13__R3_BUF_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y14__R0_BUF_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R0_INV_0 (.A(tie_lo_T19Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y14__R1_BUF_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R1_INV_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R2_INV_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y14__R2_INV_1 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y14__R3_BUF_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y15__R0_BUF_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R0_INV_0 (.A(tie_lo_T19Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y15__R1_BUF_0 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R1_INV_0 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R2_INV_0 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y15__R2_INV_1 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y15__R3_BUF_0 (.A(tie_lo_T19Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y16__R0_BUF_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R0_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y16__R1_BUF_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R1_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R2_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y16__R2_INV_1 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y16__R3_BUF_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y17__R0_BUF_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R0_INV_0 (.A(tie_lo_T19Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y17__R1_BUF_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R1_INV_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R2_INV_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y17__R2_INV_1 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y17__R3_BUF_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y18__R0_BUF_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R0_INV_0 (.A(tie_lo_T19Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y18__R1_BUF_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R1_INV_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R2_INV_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y18__R2_INV_1 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y18__R3_BUF_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y19__R0_BUF_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R0_INV_0 (.A(tie_lo_T19Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y19__R1_BUF_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R1_INV_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R2_INV_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y19__R2_INV_1 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y19__R3_BUF_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y1__R0_BUF_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R0_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y1__R1_BUF_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R1_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R2_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y1__R2_INV_1 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y1__R3_BUF_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y20__R0_BUF_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R0_INV_0 (.A(tie_lo_T19Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y20__R1_BUF_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R1_INV_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R2_INV_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y20__R2_INV_1 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y20__R3_BUF_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y21__R0_BUF_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R0_INV_0 (.A(tie_lo_T19Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y21__R1_BUF_0 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R1_INV_0 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R2_INV_0 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y21__R2_INV_1 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y21__R3_BUF_0 (.A(tie_lo_T19Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y22__R0_BUF_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R0_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y22__R1_BUF_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R1_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R2_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y22__R2_INV_1 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y22__R3_BUF_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y23__R0_BUF_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R0_INV_0 (.A(tie_lo_T19Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y23__R1_BUF_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R1_INV_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R2_INV_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y23__R2_INV_1 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y23__R3_BUF_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y24__R0_BUF_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R0_INV_0 (.A(tie_lo_T19Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y24__R1_BUF_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R1_INV_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R2_INV_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y24__R2_INV_1 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y24__R3_BUF_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y25__R0_BUF_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R0_INV_0 (.A(tie_lo_T19Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y25__R1_BUF_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R1_INV_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R2_INV_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y25__R2_INV_1 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y25__R3_BUF_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y26__R0_BUF_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R0_INV_0 (.A(tie_lo_T19Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y26__R1_BUF_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R1_INV_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R2_INV_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y26__R2_INV_1 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y26__R3_BUF_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y27__R0_BUF_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R0_INV_0 (.A(tie_lo_T19Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y27__R1_BUF_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R1_INV_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R2_INV_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y27__R2_INV_1 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y27__R3_BUF_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y28__R0_BUF_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R0_INV_0 (.A(tie_lo_T19Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y28__R1_BUF_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R1_INV_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R2_INV_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y28__R2_INV_1 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y28__R3_BUF_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y29__R0_BUF_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R0_INV_0 (.A(tie_lo_T19Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y29__R1_BUF_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R1_INV_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R2_INV_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y29__R2_INV_1 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y29__R3_BUF_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y2__R0_BUF_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R0_INV_0 (.A(tie_lo_T19Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y2__R1_BUF_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R1_INV_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R2_INV_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y2__R2_INV_1 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y2__R3_BUF_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y30__R0_BUF_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R0_INV_0 (.A(tie_lo_T19Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y30__R1_BUF_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R1_INV_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R2_INV_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y30__R2_INV_1 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y30__R3_BUF_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y31__R0_BUF_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R0_INV_0 (.A(tie_lo_T19Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y31__R1_BUF_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R1_INV_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R2_INV_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y31__R2_INV_1 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y31__R3_BUF_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y32__R0_BUF_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R0_INV_0 (.A(tie_lo_T19Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y32__R1_BUF_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R1_INV_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R2_INV_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y32__R2_INV_1 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y32__R3_BUF_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y33__R0_BUF_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R0_INV_0 (.A(tie_lo_T19Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y33__R1_BUF_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R1_INV_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R2_INV_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y33__R2_INV_1 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y33__R3_BUF_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y34__R0_BUF_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R0_INV_0 (.A(tie_lo_T19Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y34__R1_BUF_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R1_INV_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R2_INV_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y34__R2_INV_1 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y34__R3_BUF_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y35__R0_BUF_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R0_INV_0 (.A(tie_lo_T19Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y35__R1_BUF_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R1_INV_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R2_INV_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y35__R2_INV_1 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y35__R3_BUF_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y36__R0_BUF_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R0_INV_0 (.A(tie_lo_T19Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y36__R1_BUF_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R1_INV_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R2_INV_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y36__R2_INV_1 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y36__R3_BUF_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y37__R0_BUF_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R0_INV_0 (.A(tie_lo_T19Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y37__R1_BUF_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R1_INV_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R2_INV_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y37__R2_INV_1 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y37__R3_BUF_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y38__R0_BUF_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R0_INV_0 (.A(tie_lo_T19Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y38__R1_BUF_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R1_INV_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R2_INV_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y38__R2_INV_1 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y38__R3_BUF_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y39__R0_BUF_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R0_INV_0 (.A(tie_lo_T19Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y39__R1_BUF_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R1_INV_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R2_INV_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y39__R2_INV_1 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y39__R3_BUF_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y3__R0_BUF_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R0_INV_0 (.A(tie_lo_T19Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y3__R1_BUF_0 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R1_INV_0 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R2_INV_0 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y3__R2_INV_1 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y3__R3_BUF_0 (.A(tie_lo_T19Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y40__R0_BUF_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R0_INV_0 (.A(tie_lo_T19Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y40__R1_BUF_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R1_INV_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R2_INV_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y40__R2_INV_1 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y40__R3_BUF_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y41__R0_BUF_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R0_INV_0 (.A(tie_lo_T19Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y41__R1_BUF_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R1_INV_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R2_INV_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y41__R2_INV_1 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y41__R3_BUF_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y42__R0_BUF_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R0_INV_0 (.A(tie_lo_T19Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y42__R1_BUF_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R1_INV_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R2_INV_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y42__R2_INV_1 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y42__R3_BUF_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y43__R0_BUF_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R0_INV_0 (.A(tie_lo_T19Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y43__R1_BUF_0 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R1_INV_0 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R2_INV_0 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y43__R2_INV_1 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y43__R3_BUF_0 (.A(tie_lo_T19Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y44__R0_BUF_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R0_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y44__R1_BUF_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R1_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R2_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y44__R2_INV_1 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y44__R3_BUF_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y45__R0_BUF_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R0_INV_0 (.A(tie_lo_T19Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y45__R1_BUF_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R1_INV_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R2_INV_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y45__R2_INV_1 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y45__R3_BUF_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y46__R0_BUF_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R0_INV_0 (.A(tie_lo_T19Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y46__R1_BUF_0 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R1_INV_0 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R2_INV_0 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y46__R2_INV_1 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y46__R3_BUF_0 (.A(tie_lo_T19Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y47__R0_BUF_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R0_INV_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y47__R1_BUF_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R1_INV_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R2_INV_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y47__R2_INV_1 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y47__R3_BUF_0 (.A(tie_lo_T19Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y48__R0_BUF_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R0_INV_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y48__R1_BUF_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R1_INV_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R2_INV_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y48__R2_INV_1 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y48__R3_BUF_0 (.A(tie_lo_T19Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y49__R0_BUF_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R0_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y49__R1_BUF_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R1_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R2_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y49__R2_INV_1 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y49__R3_BUF_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y4__R0_BUF_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R0_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y4__R1_BUF_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R1_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R2_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y4__R2_INV_1 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y4__R3_BUF_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y50__R0_BUF_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R0_INV_0 (.A(tie_lo_T19Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y50__R1_BUF_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R1_INV_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R2_INV_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y50__R2_INV_1 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y50__R3_BUF_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y51__R0_BUF_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R0_INV_0 (.A(tie_lo_T19Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y51__R1_BUF_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R1_INV_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R2_INV_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y51__R2_INV_1 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y51__R3_BUF_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y52__R0_BUF_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R0_INV_0 (.A(tie_lo_T19Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y52__R1_BUF_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R1_INV_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R2_INV_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y52__R2_INV_1 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y52__R3_BUF_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y53__R0_BUF_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R0_INV_0 (.A(tie_lo_T19Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y53__R1_BUF_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R1_INV_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R2_INV_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y53__R2_INV_1 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y53__R3_BUF_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y54__R0_BUF_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R0_INV_0 (.A(tie_lo_T19Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y54__R1_BUF_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R1_INV_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R2_INV_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y54__R2_INV_1 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y54__R3_BUF_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y55__R0_BUF_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R0_INV_0 (.A(tie_lo_T19Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y55__R1_BUF_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R1_INV_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R2_INV_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y55__R2_INV_1 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y55__R3_BUF_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y56__R0_BUF_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R0_INV_0 (.A(tie_lo_T19Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y56__R1_BUF_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R1_INV_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R2_INV_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y56__R2_INV_1 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y56__R3_BUF_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y57__R0_BUF_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R0_INV_0 (.A(tie_lo_T19Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y57__R1_BUF_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R1_INV_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R2_INV_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y57__R2_INV_1 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y57__R3_BUF_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y58__R0_BUF_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R0_INV_0 (.A(tie_lo_T19Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y58__R1_BUF_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R1_INV_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R2_INV_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y58__R2_INV_1 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y58__R3_BUF_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y59__R0_BUF_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R0_INV_0 (.A(tie_lo_T19Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y59__R1_BUF_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R1_INV_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R2_INV_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y59__R2_INV_1 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y59__R3_BUF_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y5__R0_BUF_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R0_INV_0 (.A(tie_lo_T19Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y5__R1_BUF_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R1_INV_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R2_INV_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y5__R2_INV_1 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y5__R3_BUF_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y60__R0_BUF_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R0_INV_0 (.A(tie_lo_T19Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y60__R1_BUF_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R1_INV_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R2_INV_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y60__R2_INV_1 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y60__R3_BUF_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y61__R0_BUF_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R0_INV_0 (.A(tie_lo_T19Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y61__R1_BUF_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R1_INV_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R2_INV_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y61__R2_INV_1 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y61__R3_BUF_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y62__R0_BUF_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R0_INV_0 (.A(tie_lo_T19Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y62__R1_BUF_0 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R1_INV_0 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R2_INV_0 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y62__R2_INV_1 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y62__R3_BUF_0 (.A(tie_lo_T19Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y63__R0_BUF_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R0_INV_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y63__R1_BUF_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R1_INV_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R2_INV_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y63__R2_INV_1 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y63__R3_BUF_0 (.A(tie_lo_T19Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y64__R0_BUF_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R0_INV_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y64__R1_BUF_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R1_INV_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R2_INV_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y64__R2_INV_1 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y64__R3_BUF_0 (.A(tie_lo_T19Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y65__R0_BUF_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R0_INV_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y65__R1_BUF_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R1_INV_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R2_INV_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y65__R2_INV_1 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y65__R3_BUF_0 (.A(tie_lo_T19Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y66__R0_BUF_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R0_INV_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y66__R1_BUF_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R1_INV_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R2_INV_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y66__R2_INV_1 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y66__R3_BUF_0 (.A(tie_lo_T19Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y67__R0_BUF_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R0_INV_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y67__R1_BUF_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R1_INV_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R2_INV_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y67__R2_INV_1 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y67__R3_BUF_0 (.A(tie_lo_T19Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y68__R0_BUF_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R0_INV_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y68__R1_BUF_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R1_INV_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R2_INV_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y68__R2_INV_1 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y68__R3_BUF_0 (.A(tie_lo_T19Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y69__R0_BUF_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R0_INV_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y69__R1_BUF_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R1_INV_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R2_INV_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y69__R2_INV_1 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y69__R3_BUF_0 (.A(tie_lo_T19Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y6__R0_BUF_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R0_INV_0 (.A(tie_lo_T19Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y6__R1_BUF_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R1_INV_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R2_INV_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y6__R2_INV_1 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y6__R3_BUF_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y70__R0_BUF_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R0_INV_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y70__R1_BUF_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R1_INV_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R2_INV_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y70__R2_INV_1 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y70__R3_BUF_0 (.A(tie_lo_T19Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y71__R0_BUF_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R0_INV_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y71__R1_BUF_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R1_INV_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R2_INV_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y71__R2_INV_1 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y71__R3_BUF_0 (.A(tie_lo_T19Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y72__R0_BUF_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R0_INV_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y72__R1_BUF_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R1_INV_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R2_INV_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y72__R2_INV_1 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y72__R3_BUF_0 (.A(tie_lo_T19Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y73__R0_BUF_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R0_INV_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y73__R1_BUF_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R1_INV_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R2_INV_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y73__R2_INV_1 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y73__R3_BUF_0 (.A(tie_lo_T19Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y74__R0_BUF_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R0_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y74__R1_BUF_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R1_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R2_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y74__R2_INV_1 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y74__R3_BUF_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y75__R0_BUF_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R0_INV_0 (.A(tie_lo_T19Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y75__R1_BUF_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R1_INV_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R2_INV_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y75__R2_INV_1 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y75__R3_BUF_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y76__R0_BUF_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R0_INV_0 (.A(tie_lo_T19Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y76__R1_BUF_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R1_INV_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R2_INV_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y76__R2_INV_1 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y76__R3_BUF_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y77__R0_BUF_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R0_INV_0 (.A(tie_lo_T19Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y77__R1_BUF_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R1_INV_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R2_INV_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y77__R2_INV_1 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y77__R3_BUF_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y78__R0_BUF_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R0_INV_0 (.A(tie_lo_T19Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y78__R1_BUF_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R1_INV_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R2_INV_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y78__R2_INV_1 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y78__R3_BUF_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y79__R0_BUF_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R0_INV_0 (.A(tie_lo_T19Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y79__R1_BUF_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R1_INV_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R2_INV_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y79__R2_INV_1 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y79__R3_BUF_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y7__R0_BUF_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R0_INV_0 (.A(tie_lo_T19Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y7__R1_BUF_0 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R1_INV_0 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R2_INV_0 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y7__R2_INV_1 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y7__R3_BUF_0 (.A(tie_lo_T19Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y80__R0_BUF_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R0_INV_0 (.A(tie_lo_T19Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y80__R1_BUF_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R1_INV_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R2_INV_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y80__R2_INV_1 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y80__R3_BUF_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y81__R0_BUF_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R0_INV_0 (.A(tie_lo_T19Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y81__R1_BUF_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R1_INV_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R2_INV_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y81__R2_INV_1 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y81__R3_BUF_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y82__R0_BUF_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R0_INV_0 (.A(tie_lo_T19Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y82__R1_BUF_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R1_INV_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R2_INV_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y82__R2_INV_1 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y82__R3_BUF_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y83__R0_BUF_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R0_INV_0 (.A(tie_lo_T19Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y83__R1_BUF_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R1_INV_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R2_INV_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y83__R2_INV_1 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y83__R3_BUF_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y84__R0_BUF_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R0_INV_0 (.A(tie_lo_T19Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y84__R1_BUF_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R1_INV_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R2_INV_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y84__R2_INV_1 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y84__R3_BUF_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y85__R0_BUF_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R0_INV_0 (.A(tie_lo_T19Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y85__R1_BUF_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R1_INV_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R2_INV_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y85__R2_INV_1 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y85__R3_BUF_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y86__R0_BUF_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R0_INV_0 (.A(tie_lo_T19Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y86__R1_BUF_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R1_INV_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R2_INV_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y86__R2_INV_1 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y86__R3_BUF_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y87__R0_BUF_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R0_INV_0 (.A(tie_lo_T19Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y87__R1_BUF_0 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R1_INV_0 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R2_INV_0 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y87__R2_INV_1 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y87__R3_BUF_0 (.A(tie_lo_T19Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y88__R0_BUF_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R0_INV_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y88__R1_BUF_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R1_INV_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R2_INV_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y88__R2_INV_1 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y88__R3_BUF_0 (.A(tie_lo_T19Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y89__R0_BUF_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R0_INV_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y89__R1_BUF_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R1_INV_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R2_INV_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y89__R2_INV_1 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y89__R3_BUF_0 (.A(tie_lo_T19Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y8__R0_BUF_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R0_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y8__R1_BUF_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R1_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R2_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y8__R2_INV_1 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y8__R3_BUF_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y9__R0_BUF_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R0_INV_0 (.A(tie_lo_T19Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y9__R1_BUF_0 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R1_INV_0 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T19Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R2_INV_0 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T19Y9__R2_INV_1 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T19Y9__R3_BUF_0 (.A(tie_lo_T19Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y0__R0_BUF_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R0_INV_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y0__R1_BUF_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R1_INV_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R2_INV_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y0__R2_INV_1 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y0__R3_BUF_0 (.A(tie_lo_T1Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y10__R0_BUF_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R0_INV_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y10__R1_BUF_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R1_INV_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R2_INV_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y10__R2_INV_1 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y10__R3_BUF_0 (.A(tie_lo_T1Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y11__R0_BUF_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R0_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y11__R1_BUF_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R1_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R2_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y11__R2_INV_1 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y11__R3_BUF_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y12__R0_BUF_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R0_INV_0 (.A(tie_lo_T1Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y12__R1_BUF_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R1_INV_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R2_INV_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y12__R2_INV_1 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y12__R3_BUF_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y13__R0_BUF_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R0_INV_0 (.A(tie_lo_T1Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y13__R1_BUF_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R1_INV_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R2_INV_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y13__R2_INV_1 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y13__R3_BUF_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y14__R0_BUF_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R0_INV_0 (.A(tie_lo_T1Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y14__R1_BUF_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R1_INV_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R2_INV_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y14__R2_INV_1 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y14__R3_BUF_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y15__R0_BUF_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R0_INV_0 (.A(tie_lo_T1Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y15__R1_BUF_0 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R1_INV_0 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R2_INV_0 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y15__R2_INV_1 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y15__R3_BUF_0 (.A(tie_lo_T1Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y16__R0_BUF_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R0_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y16__R1_BUF_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R1_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R2_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y16__R2_INV_1 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y16__R3_BUF_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y17__R0_BUF_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R0_INV_0 (.A(tie_lo_T1Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y17__R1_BUF_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R1_INV_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R2_INV_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y17__R2_INV_1 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y17__R3_BUF_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y18__R0_BUF_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R0_INV_0 (.A(tie_lo_T1Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y18__R1_BUF_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R1_INV_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R2_INV_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y18__R2_INV_1 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y18__R3_BUF_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y19__R0_BUF_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R0_INV_0 (.A(tie_lo_T1Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y19__R1_BUF_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R1_INV_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R2_INV_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y19__R2_INV_1 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y19__R3_BUF_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y1__R0_BUF_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R0_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y1__R1_BUF_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R1_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R2_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y1__R2_INV_1 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y1__R3_BUF_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y20__R0_BUF_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R0_INV_0 (.A(tie_lo_T1Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y20__R1_BUF_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R1_INV_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R2_INV_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y20__R2_INV_1 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y20__R3_BUF_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y21__R0_BUF_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R0_INV_0 (.A(tie_lo_T1Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y21__R1_BUF_0 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R1_INV_0 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R2_INV_0 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y21__R2_INV_1 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y21__R3_BUF_0 (.A(tie_lo_T1Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y22__R0_BUF_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R0_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y22__R1_BUF_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R1_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R2_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y22__R2_INV_1 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y22__R3_BUF_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y23__R0_BUF_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R0_INV_0 (.A(tie_lo_T1Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y23__R1_BUF_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R1_INV_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R2_INV_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y23__R2_INV_1 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y23__R3_BUF_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y24__R0_BUF_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R0_INV_0 (.A(tie_lo_T1Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y24__R1_BUF_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R1_INV_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R2_INV_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y24__R2_INV_1 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y24__R3_BUF_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y25__R0_BUF_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R0_INV_0 (.A(tie_lo_T1Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y25__R1_BUF_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R1_INV_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R2_INV_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y25__R2_INV_1 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y25__R3_BUF_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y26__R0_BUF_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R0_INV_0 (.A(tie_lo_T1Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y26__R1_BUF_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R1_INV_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R2_INV_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y26__R2_INV_1 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y26__R3_BUF_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y27__R0_BUF_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R0_INV_0 (.A(tie_lo_T1Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y27__R1_BUF_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R1_INV_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R2_INV_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y27__R2_INV_1 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y27__R3_BUF_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y28__R0_BUF_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R0_INV_0 (.A(tie_lo_T1Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y28__R1_BUF_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R1_INV_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R2_INV_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y28__R2_INV_1 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y28__R3_BUF_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y29__R0_BUF_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R0_INV_0 (.A(tie_lo_T1Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y29__R1_BUF_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R1_INV_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R2_INV_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y29__R2_INV_1 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y29__R3_BUF_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y2__R0_BUF_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R0_INV_0 (.A(tie_lo_T1Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y2__R1_BUF_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R1_INV_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R2_INV_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y2__R2_INV_1 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y2__R3_BUF_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y30__R0_BUF_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R0_INV_0 (.A(tie_lo_T1Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y30__R1_BUF_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R1_INV_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R2_INV_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y30__R2_INV_1 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y30__R3_BUF_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y31__R0_BUF_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R0_INV_0 (.A(tie_lo_T1Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y31__R1_BUF_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R1_INV_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R2_INV_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y31__R2_INV_1 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y31__R3_BUF_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y32__R0_BUF_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R0_INV_0 (.A(tie_lo_T1Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y32__R1_BUF_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R1_INV_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R2_INV_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y32__R2_INV_1 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y32__R3_BUF_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y33__R0_BUF_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R0_INV_0 (.A(tie_lo_T1Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y33__R1_BUF_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R1_INV_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R2_INV_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y33__R2_INV_1 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y33__R3_BUF_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y34__R0_BUF_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R0_INV_0 (.A(tie_lo_T1Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y34__R1_BUF_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R1_INV_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R2_INV_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y34__R2_INV_1 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y34__R3_BUF_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y35__R0_BUF_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R0_INV_0 (.A(tie_lo_T1Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y35__R1_BUF_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R1_INV_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R2_INV_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y35__R2_INV_1 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y35__R3_BUF_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y36__R0_BUF_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R0_INV_0 (.A(tie_lo_T1Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y36__R1_BUF_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R1_INV_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R2_INV_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y36__R2_INV_1 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y36__R3_BUF_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y37__R0_BUF_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R0_INV_0 (.A(tie_lo_T1Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y37__R1_BUF_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R1_INV_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R2_INV_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y37__R2_INV_1 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y37__R3_BUF_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y38__R0_BUF_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R0_INV_0 (.A(tie_lo_T1Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y38__R1_BUF_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R1_INV_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R2_INV_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y38__R2_INV_1 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y38__R3_BUF_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y39__R0_BUF_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R0_INV_0 (.A(tie_lo_T1Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y39__R1_BUF_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R1_INV_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R2_INV_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y39__R2_INV_1 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y39__R3_BUF_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y3__R0_BUF_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R0_INV_0 (.A(tie_lo_T1Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y3__R1_BUF_0 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R1_INV_0 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R2_INV_0 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y3__R2_INV_1 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y3__R3_BUF_0 (.A(tie_lo_T1Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y40__R0_BUF_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R0_INV_0 (.A(tie_lo_T1Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y40__R1_BUF_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R1_INV_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R2_INV_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y40__R2_INV_1 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y40__R3_BUF_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y41__R0_BUF_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R0_INV_0 (.A(tie_lo_T1Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y41__R1_BUF_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R1_INV_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R2_INV_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y41__R2_INV_1 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y41__R3_BUF_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y42__R0_BUF_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R0_INV_0 (.A(tie_lo_T1Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y42__R1_BUF_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R1_INV_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R2_INV_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y42__R2_INV_1 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y42__R3_BUF_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y43__R0_BUF_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R0_INV_0 (.A(tie_lo_T1Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y43__R1_BUF_0 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R1_INV_0 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R2_INV_0 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y43__R2_INV_1 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y43__R3_BUF_0 (.A(tie_lo_T1Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y44__R0_BUF_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R0_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y44__R1_BUF_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R1_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R2_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y44__R2_INV_1 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y44__R3_BUF_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y45__R0_BUF_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R0_INV_0 (.A(tie_lo_T1Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y45__R1_BUF_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R1_INV_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R2_INV_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y45__R2_INV_1 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y45__R3_BUF_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y46__R0_BUF_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R0_INV_0 (.A(tie_lo_T1Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y46__R1_BUF_0 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R1_INV_0 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R2_INV_0 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y46__R2_INV_1 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y46__R3_BUF_0 (.A(tie_lo_T1Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y47__R0_BUF_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R0_INV_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y47__R1_BUF_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R1_INV_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R2_INV_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y47__R2_INV_1 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y47__R3_BUF_0 (.A(tie_lo_T1Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y48__R0_BUF_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R0_INV_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y48__R1_BUF_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R1_INV_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R2_INV_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y48__R2_INV_1 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y48__R3_BUF_0 (.A(tie_lo_T1Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y49__R0_BUF_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R0_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y49__R1_BUF_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R1_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R2_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y49__R2_INV_1 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y49__R3_BUF_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y4__R0_BUF_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R0_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y4__R1_BUF_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R1_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R2_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y4__R2_INV_1 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y4__R3_BUF_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y50__R0_BUF_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R0_INV_0 (.A(tie_lo_T1Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y50__R1_BUF_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R1_INV_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R2_INV_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y50__R2_INV_1 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y50__R3_BUF_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y51__R0_BUF_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R0_INV_0 (.A(tie_lo_T1Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y51__R1_BUF_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R1_INV_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R2_INV_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y51__R2_INV_1 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y51__R3_BUF_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y52__R0_BUF_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R0_INV_0 (.A(tie_lo_T1Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y52__R1_BUF_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R1_INV_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R2_INV_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y52__R2_INV_1 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y52__R3_BUF_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y53__R0_BUF_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R0_INV_0 (.A(tie_lo_T1Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y53__R1_BUF_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R1_INV_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R2_INV_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y53__R2_INV_1 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y53__R3_BUF_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y54__R0_BUF_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R0_INV_0 (.A(tie_lo_T1Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y54__R1_BUF_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R1_INV_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R2_INV_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y54__R2_INV_1 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y54__R3_BUF_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y55__R0_BUF_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R0_INV_0 (.A(tie_lo_T1Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y55__R1_BUF_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R1_INV_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R2_INV_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y55__R2_INV_1 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y55__R3_BUF_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y56__R0_BUF_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R0_INV_0 (.A(tie_lo_T1Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y56__R1_BUF_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R1_INV_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R2_INV_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y56__R2_INV_1 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y56__R3_BUF_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y57__R0_BUF_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R0_INV_0 (.A(tie_lo_T1Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y57__R1_BUF_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R1_INV_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R2_INV_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y57__R2_INV_1 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y57__R3_BUF_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y58__R0_BUF_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R0_INV_0 (.A(tie_lo_T1Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y58__R1_BUF_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R1_INV_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R2_INV_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y58__R2_INV_1 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y58__R3_BUF_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y59__R0_BUF_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R0_INV_0 (.A(tie_lo_T1Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y59__R1_BUF_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R1_INV_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R2_INV_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y59__R2_INV_1 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y59__R3_BUF_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y5__R0_BUF_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R0_INV_0 (.A(tie_lo_T1Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y5__R1_BUF_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R1_INV_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R2_INV_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y5__R2_INV_1 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y5__R3_BUF_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y60__R0_BUF_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R0_INV_0 (.A(tie_lo_T1Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y60__R1_BUF_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R1_INV_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R2_INV_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y60__R2_INV_1 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y60__R3_BUF_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y61__R0_BUF_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R0_INV_0 (.A(tie_lo_T1Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y61__R1_BUF_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R1_INV_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R2_INV_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y61__R2_INV_1 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y61__R3_BUF_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y62__R0_BUF_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R0_INV_0 (.A(tie_lo_T1Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y62__R1_BUF_0 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R1_INV_0 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R2_INV_0 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y62__R2_INV_1 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y62__R3_BUF_0 (.A(tie_lo_T1Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y63__R0_BUF_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R0_INV_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y63__R1_BUF_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R1_INV_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R2_INV_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y63__R2_INV_1 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y63__R3_BUF_0 (.A(tie_lo_T1Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y64__R0_BUF_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R0_INV_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y64__R1_BUF_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R1_INV_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R2_INV_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y64__R2_INV_1 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y64__R3_BUF_0 (.A(tie_lo_T1Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y65__R0_BUF_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R0_INV_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y65__R1_BUF_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R1_INV_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R2_INV_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y65__R2_INV_1 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y65__R3_BUF_0 (.A(tie_lo_T1Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y66__R0_BUF_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R0_INV_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y66__R1_BUF_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R1_INV_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R2_INV_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y66__R2_INV_1 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y66__R3_BUF_0 (.A(tie_lo_T1Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y67__R0_BUF_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R0_INV_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y67__R1_BUF_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R1_INV_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R2_INV_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y67__R2_INV_1 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y67__R3_BUF_0 (.A(tie_lo_T1Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y68__R0_BUF_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R0_INV_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y68__R1_BUF_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R1_INV_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R2_INV_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y68__R2_INV_1 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y68__R3_BUF_0 (.A(tie_lo_T1Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y69__R0_BUF_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R0_INV_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y69__R1_BUF_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R1_INV_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R2_INV_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y69__R2_INV_1 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y69__R3_BUF_0 (.A(tie_lo_T1Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y6__R0_BUF_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R0_INV_0 (.A(tie_lo_T1Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y6__R1_BUF_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R1_INV_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R2_INV_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y6__R2_INV_1 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y6__R3_BUF_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y70__R0_BUF_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R0_INV_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y70__R1_BUF_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R1_INV_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R2_INV_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y70__R2_INV_1 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y70__R3_BUF_0 (.A(tie_lo_T1Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y71__R0_BUF_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R0_INV_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y71__R1_BUF_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R1_INV_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R2_INV_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y71__R2_INV_1 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y71__R3_BUF_0 (.A(tie_lo_T1Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y72__R0_BUF_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R0_INV_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y72__R1_BUF_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R1_INV_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R2_INV_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y72__R2_INV_1 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y72__R3_BUF_0 (.A(tie_lo_T1Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y73__R0_BUF_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R0_INV_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y73__R1_BUF_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R1_INV_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R2_INV_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y73__R2_INV_1 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y73__R3_BUF_0 (.A(tie_lo_T1Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y74__R0_BUF_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R0_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y74__R1_BUF_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R1_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R2_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y74__R2_INV_1 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y74__R3_BUF_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y75__R0_BUF_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R0_INV_0 (.A(tie_lo_T1Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y75__R1_BUF_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R1_INV_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R2_INV_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y75__R2_INV_1 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y75__R3_BUF_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y76__R0_BUF_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R0_INV_0 (.A(tie_lo_T1Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y76__R1_BUF_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R1_INV_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R2_INV_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y76__R2_INV_1 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y76__R3_BUF_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y77__R0_BUF_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R0_INV_0 (.A(tie_lo_T1Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y77__R1_BUF_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R1_INV_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R2_INV_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y77__R2_INV_1 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y77__R3_BUF_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y78__R0_BUF_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R0_INV_0 (.A(tie_lo_T1Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y78__R1_BUF_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R1_INV_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R2_INV_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y78__R2_INV_1 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y78__R3_BUF_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y79__R0_BUF_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R0_INV_0 (.A(tie_lo_T1Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y79__R1_BUF_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R1_INV_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R2_INV_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y79__R2_INV_1 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y79__R3_BUF_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y7__R0_BUF_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R0_INV_0 (.A(tie_lo_T1Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y7__R1_BUF_0 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R1_INV_0 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R2_INV_0 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y7__R2_INV_1 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y7__R3_BUF_0 (.A(tie_lo_T1Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y80__R0_BUF_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R0_INV_0 (.A(tie_lo_T1Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y80__R1_BUF_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R1_INV_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R2_INV_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y80__R2_INV_1 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y80__R3_BUF_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y81__R0_BUF_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R0_INV_0 (.A(tie_lo_T1Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y81__R1_BUF_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R1_INV_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R2_INV_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y81__R2_INV_1 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y81__R3_BUF_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y82__R0_BUF_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R0_INV_0 (.A(tie_lo_T1Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y82__R1_BUF_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R1_INV_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R2_INV_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y82__R2_INV_1 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y82__R3_BUF_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y83__R0_BUF_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R0_INV_0 (.A(tie_lo_T1Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y83__R1_BUF_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R1_INV_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R2_INV_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y83__R2_INV_1 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y83__R3_BUF_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y84__R0_BUF_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R0_INV_0 (.A(tie_lo_T1Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y84__R1_BUF_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R1_INV_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R2_INV_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y84__R2_INV_1 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y84__R3_BUF_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y85__R0_BUF_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R0_INV_0 (.A(tie_lo_T1Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y85__R1_BUF_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R1_INV_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R2_INV_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y85__R2_INV_1 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y85__R3_BUF_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y86__R0_BUF_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R0_INV_0 (.A(tie_lo_T1Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y86__R1_BUF_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R1_INV_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R2_INV_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y86__R2_INV_1 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y86__R3_BUF_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y87__R0_BUF_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R0_INV_0 (.A(tie_lo_T1Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y87__R1_BUF_0 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R1_INV_0 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R2_INV_0 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y87__R2_INV_1 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y87__R3_BUF_0 (.A(tie_lo_T1Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y88__R0_BUF_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R0_INV_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y88__R1_BUF_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R1_INV_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R2_INV_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y88__R2_INV_1 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y88__R3_BUF_0 (.A(tie_lo_T1Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y89__R0_BUF_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R0_INV_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y89__R1_BUF_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R1_INV_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R2_INV_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y89__R2_INV_1 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y89__R3_BUF_0 (.A(tie_lo_T1Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y8__R0_BUF_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R0_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y8__R1_BUF_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R1_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R2_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y8__R2_INV_1 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y8__R3_BUF_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y9__R0_BUF_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R0_INV_0 (.A(tie_lo_T1Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y9__R1_BUF_0 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R1_INV_0 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T1Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R2_INV_0 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T1Y9__R2_INV_1 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T1Y9__R3_BUF_0 (.A(tie_lo_T1Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y0__R0_BUF_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R0_INV_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y0__R1_BUF_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R1_INV_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R2_INV_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y0__R2_INV_1 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y0__R3_BUF_0 (.A(tie_lo_T20Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y10__R0_BUF_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R0_INV_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y10__R1_BUF_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R1_INV_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R2_INV_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y10__R2_INV_1 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y10__R3_BUF_0 (.A(tie_lo_T20Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y11__R0_BUF_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R0_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y11__R1_BUF_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R1_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R2_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y11__R2_INV_1 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y11__R3_BUF_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y12__R0_BUF_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R0_INV_0 (.A(tie_lo_T20Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y12__R1_BUF_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R1_INV_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R2_INV_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y12__R2_INV_1 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y12__R3_BUF_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y13__R0_BUF_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R0_INV_0 (.A(tie_lo_T20Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y13__R1_BUF_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R1_INV_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R2_INV_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y13__R2_INV_1 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y13__R3_BUF_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y14__R0_BUF_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R0_INV_0 (.A(tie_lo_T20Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y14__R1_BUF_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R1_INV_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R2_INV_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y14__R2_INV_1 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y14__R3_BUF_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y15__R0_BUF_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R0_INV_0 (.A(tie_lo_T20Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y15__R1_BUF_0 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R1_INV_0 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R2_INV_0 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y15__R2_INV_1 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y15__R3_BUF_0 (.A(tie_lo_T20Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y16__R0_BUF_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R0_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y16__R1_BUF_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R1_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R2_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y16__R2_INV_1 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y16__R3_BUF_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y17__R0_BUF_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R0_INV_0 (.A(tie_lo_T20Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y17__R1_BUF_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R1_INV_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R2_INV_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y17__R2_INV_1 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y17__R3_BUF_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y18__R0_BUF_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R0_INV_0 (.A(tie_lo_T20Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y18__R1_BUF_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R1_INV_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R2_INV_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y18__R2_INV_1 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y18__R3_BUF_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y19__R0_BUF_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R0_INV_0 (.A(tie_lo_T20Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y19__R1_BUF_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R1_INV_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R2_INV_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y19__R2_INV_1 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y19__R3_BUF_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y1__R0_BUF_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R0_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y1__R1_BUF_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R1_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R2_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y1__R2_INV_1 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y1__R3_BUF_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y20__R0_BUF_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R0_INV_0 (.A(tie_lo_T20Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y20__R1_BUF_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R1_INV_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R2_INV_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y20__R2_INV_1 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y20__R3_BUF_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y21__R0_BUF_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R0_INV_0 (.A(tie_lo_T20Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y21__R1_BUF_0 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R1_INV_0 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R2_INV_0 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y21__R2_INV_1 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y21__R3_BUF_0 (.A(tie_lo_T20Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y22__R0_BUF_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R0_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y22__R1_BUF_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R1_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R2_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y22__R2_INV_1 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y22__R3_BUF_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y23__R0_BUF_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R0_INV_0 (.A(tie_lo_T20Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y23__R1_BUF_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R1_INV_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R2_INV_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y23__R2_INV_1 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y23__R3_BUF_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y24__R0_BUF_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R0_INV_0 (.A(tie_lo_T20Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y24__R1_BUF_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R1_INV_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R2_INV_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y24__R2_INV_1 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y24__R3_BUF_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y25__R0_BUF_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R0_INV_0 (.A(tie_lo_T20Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y25__R1_BUF_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R1_INV_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R2_INV_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y25__R2_INV_1 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y25__R3_BUF_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y26__R0_BUF_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R0_INV_0 (.A(tie_lo_T20Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y26__R1_BUF_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R1_INV_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R2_INV_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y26__R2_INV_1 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y26__R3_BUF_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y27__R0_BUF_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R0_INV_0 (.A(tie_lo_T20Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y27__R1_BUF_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R1_INV_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R2_INV_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y27__R2_INV_1 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y27__R3_BUF_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y28__R0_BUF_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R0_INV_0 (.A(tie_lo_T20Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y28__R1_BUF_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R1_INV_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R2_INV_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y28__R2_INV_1 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y28__R3_BUF_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y29__R0_BUF_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R0_INV_0 (.A(tie_lo_T20Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y29__R1_BUF_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R1_INV_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R2_INV_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y29__R2_INV_1 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y29__R3_BUF_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y2__R0_BUF_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R0_INV_0 (.A(tie_lo_T20Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y2__R1_BUF_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R1_INV_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R2_INV_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y2__R2_INV_1 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y2__R3_BUF_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y30__R0_BUF_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R0_INV_0 (.A(tie_lo_T20Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y30__R1_BUF_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R1_INV_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R2_INV_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y30__R2_INV_1 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y30__R3_BUF_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y31__R0_BUF_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R0_INV_0 (.A(tie_lo_T20Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y31__R1_BUF_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R1_INV_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R2_INV_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y31__R2_INV_1 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y31__R3_BUF_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y32__R0_BUF_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R0_INV_0 (.A(tie_lo_T20Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y32__R1_BUF_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R1_INV_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R2_INV_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y32__R2_INV_1 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y32__R3_BUF_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y33__R0_BUF_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R0_INV_0 (.A(tie_lo_T20Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y33__R1_BUF_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R1_INV_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R2_INV_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y33__R2_INV_1 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y33__R3_BUF_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y34__R0_BUF_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R0_INV_0 (.A(tie_lo_T20Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y34__R1_BUF_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R1_INV_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R2_INV_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y34__R2_INV_1 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y34__R3_BUF_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y35__R0_BUF_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R0_INV_0 (.A(tie_lo_T20Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y35__R1_BUF_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R1_INV_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R2_INV_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y35__R2_INV_1 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y35__R3_BUF_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y36__R0_BUF_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R0_INV_0 (.A(tie_lo_T20Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y36__R1_BUF_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R1_INV_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R2_INV_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y36__R2_INV_1 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y36__R3_BUF_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y37__R0_BUF_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R0_INV_0 (.A(tie_lo_T20Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y37__R1_BUF_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R1_INV_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R2_INV_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y37__R2_INV_1 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y37__R3_BUF_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y38__R0_BUF_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R0_INV_0 (.A(tie_lo_T20Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y38__R1_BUF_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R1_INV_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R2_INV_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y38__R2_INV_1 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y38__R3_BUF_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y39__R0_BUF_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R0_INV_0 (.A(tie_lo_T20Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y39__R1_BUF_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R1_INV_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R2_INV_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y39__R2_INV_1 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y39__R3_BUF_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y3__R0_BUF_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R0_INV_0 (.A(tie_lo_T20Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y3__R1_BUF_0 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R1_INV_0 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R2_INV_0 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y3__R2_INV_1 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y3__R3_BUF_0 (.A(tie_lo_T20Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y40__R0_BUF_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R0_INV_0 (.A(tie_lo_T20Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y40__R1_BUF_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R1_INV_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R2_INV_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y40__R2_INV_1 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y40__R3_BUF_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y41__R0_BUF_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R0_INV_0 (.A(tie_lo_T20Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y41__R1_BUF_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R1_INV_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R2_INV_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y41__R2_INV_1 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y41__R3_BUF_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y42__R0_BUF_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R0_INV_0 (.A(tie_lo_T20Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y42__R1_BUF_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R1_INV_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R2_INV_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y42__R2_INV_1 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y42__R3_BUF_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y43__R0_BUF_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R0_INV_0 (.A(tie_lo_T20Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y43__R1_BUF_0 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R1_INV_0 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R2_INV_0 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y43__R2_INV_1 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y43__R3_BUF_0 (.A(tie_lo_T20Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y44__R0_BUF_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R0_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y44__R1_BUF_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R1_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R2_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y44__R2_INV_1 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y44__R3_BUF_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y45__R0_BUF_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R0_INV_0 (.A(tie_lo_T20Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y45__R1_BUF_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R1_INV_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R2_INV_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y45__R2_INV_1 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y45__R3_BUF_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y46__R0_BUF_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R0_INV_0 (.A(tie_lo_T20Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y46__R1_BUF_0 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R1_INV_0 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R2_INV_0 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y46__R2_INV_1 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y46__R3_BUF_0 (.A(tie_lo_T20Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y47__R0_BUF_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R0_INV_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y47__R1_BUF_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R1_INV_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R2_INV_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y47__R2_INV_1 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y47__R3_BUF_0 (.A(tie_lo_T20Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y48__R0_BUF_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R0_INV_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y48__R1_BUF_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R1_INV_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R2_INV_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y48__R2_INV_1 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y48__R3_BUF_0 (.A(tie_lo_T20Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y49__R0_BUF_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R0_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y49__R1_BUF_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R1_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R2_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y49__R2_INV_1 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y49__R3_BUF_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y4__R0_BUF_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R0_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y4__R1_BUF_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R1_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R2_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y4__R2_INV_1 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y4__R3_BUF_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y50__R0_BUF_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R0_INV_0 (.A(tie_lo_T20Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y50__R1_BUF_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R1_INV_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R2_INV_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y50__R2_INV_1 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y50__R3_BUF_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y51__R0_BUF_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R0_INV_0 (.A(tie_lo_T20Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y51__R1_BUF_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R1_INV_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R2_INV_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y51__R2_INV_1 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y51__R3_BUF_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y52__R0_BUF_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R0_INV_0 (.A(tie_lo_T20Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y52__R1_BUF_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R1_INV_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R2_INV_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y52__R2_INV_1 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y52__R3_BUF_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y53__R0_BUF_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R0_INV_0 (.A(tie_lo_T20Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y53__R1_BUF_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R1_INV_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R2_INV_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y53__R2_INV_1 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y53__R3_BUF_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y54__R0_BUF_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R0_INV_0 (.A(tie_lo_T20Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y54__R1_BUF_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R1_INV_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R2_INV_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y54__R2_INV_1 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y54__R3_BUF_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y55__R0_BUF_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R0_INV_0 (.A(tie_lo_T20Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y55__R1_BUF_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R1_INV_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R2_INV_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y55__R2_INV_1 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y55__R3_BUF_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y56__R0_BUF_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R0_INV_0 (.A(tie_lo_T20Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y56__R1_BUF_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R1_INV_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R2_INV_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y56__R2_INV_1 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y56__R3_BUF_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y57__R0_BUF_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R0_INV_0 (.A(tie_lo_T20Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y57__R1_BUF_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R1_INV_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R2_INV_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y57__R2_INV_1 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y57__R3_BUF_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y58__R0_BUF_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R0_INV_0 (.A(tie_lo_T20Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y58__R1_BUF_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R1_INV_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R2_INV_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y58__R2_INV_1 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y58__R3_BUF_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y59__R0_BUF_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R0_INV_0 (.A(tie_lo_T20Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y59__R1_BUF_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R1_INV_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R2_INV_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y59__R2_INV_1 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y59__R3_BUF_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y5__R0_BUF_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R0_INV_0 (.A(tie_lo_T20Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y5__R1_BUF_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R1_INV_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R2_INV_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y5__R2_INV_1 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y5__R3_BUF_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y60__R0_BUF_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R0_INV_0 (.A(tie_lo_T20Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y60__R1_BUF_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R1_INV_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R2_INV_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y60__R2_INV_1 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y60__R3_BUF_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y61__R0_BUF_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R0_INV_0 (.A(tie_lo_T20Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y61__R1_BUF_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R1_INV_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R2_INV_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y61__R2_INV_1 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y61__R3_BUF_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y62__R0_BUF_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R0_INV_0 (.A(tie_lo_T20Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y62__R1_BUF_0 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R1_INV_0 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R2_INV_0 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y62__R2_INV_1 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y62__R3_BUF_0 (.A(tie_lo_T20Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y63__R0_BUF_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R0_INV_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y63__R1_BUF_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R1_INV_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R2_INV_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y63__R2_INV_1 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y63__R3_BUF_0 (.A(tie_lo_T20Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y64__R0_BUF_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R0_INV_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y64__R1_BUF_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R1_INV_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R2_INV_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y64__R2_INV_1 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y64__R3_BUF_0 (.A(tie_lo_T20Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y65__R0_BUF_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R0_INV_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y65__R1_BUF_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R1_INV_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R2_INV_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y65__R2_INV_1 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y65__R3_BUF_0 (.A(tie_lo_T20Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y66__R0_BUF_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R0_INV_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y66__R1_BUF_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R1_INV_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R2_INV_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y66__R2_INV_1 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y66__R3_BUF_0 (.A(tie_lo_T20Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y67__R0_BUF_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R0_INV_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y67__R1_BUF_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R1_INV_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R2_INV_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y67__R2_INV_1 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y67__R3_BUF_0 (.A(tie_lo_T20Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y68__R0_BUF_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R0_INV_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y68__R1_BUF_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R1_INV_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R2_INV_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y68__R2_INV_1 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y68__R3_BUF_0 (.A(tie_lo_T20Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y69__R0_BUF_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R0_INV_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y69__R1_BUF_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R1_INV_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R2_INV_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y69__R2_INV_1 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y69__R3_BUF_0 (.A(tie_lo_T20Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y6__R0_BUF_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R0_INV_0 (.A(tie_lo_T20Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y6__R1_BUF_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R1_INV_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R2_INV_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y6__R2_INV_1 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y6__R3_BUF_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y70__R0_BUF_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R0_INV_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y70__R1_BUF_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R1_INV_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R2_INV_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y70__R2_INV_1 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y70__R3_BUF_0 (.A(tie_lo_T20Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y71__R0_BUF_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R0_INV_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y71__R1_BUF_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R1_INV_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R2_INV_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y71__R2_INV_1 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y71__R3_BUF_0 (.A(tie_lo_T20Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y72__R0_BUF_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R0_INV_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y72__R1_BUF_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R1_INV_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R2_INV_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y72__R2_INV_1 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y72__R3_BUF_0 (.A(tie_lo_T20Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y73__R0_BUF_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R0_INV_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y73__R1_BUF_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R1_INV_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R2_INV_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y73__R2_INV_1 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y73__R3_BUF_0 (.A(tie_lo_T20Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y74__R0_BUF_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R0_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y74__R1_BUF_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R1_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R2_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y74__R2_INV_1 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y74__R3_BUF_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y75__R0_BUF_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R0_INV_0 (.A(tie_lo_T20Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y75__R1_BUF_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R1_INV_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R2_INV_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y75__R2_INV_1 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y75__R3_BUF_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y76__R0_BUF_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R0_INV_0 (.A(tie_lo_T20Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y76__R1_BUF_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R1_INV_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R2_INV_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y76__R2_INV_1 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y76__R3_BUF_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y77__R0_BUF_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R0_INV_0 (.A(tie_lo_T20Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y77__R1_BUF_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R1_INV_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R2_INV_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y77__R2_INV_1 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y77__R3_BUF_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y78__R0_BUF_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R0_INV_0 (.A(tie_lo_T20Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y78__R1_BUF_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R1_INV_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R2_INV_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y78__R2_INV_1 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y78__R3_BUF_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y79__R0_BUF_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R0_INV_0 (.A(tie_lo_T20Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y79__R1_BUF_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R1_INV_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R2_INV_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y79__R2_INV_1 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y79__R3_BUF_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y7__R0_BUF_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R0_INV_0 (.A(tie_lo_T20Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y7__R1_BUF_0 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R1_INV_0 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R2_INV_0 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y7__R2_INV_1 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y7__R3_BUF_0 (.A(tie_lo_T20Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y80__R0_BUF_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R0_INV_0 (.A(tie_lo_T20Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y80__R1_BUF_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R1_INV_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R2_INV_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y80__R2_INV_1 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y80__R3_BUF_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y81__R0_BUF_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R0_INV_0 (.A(tie_lo_T20Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y81__R1_BUF_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R1_INV_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R2_INV_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y81__R2_INV_1 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y81__R3_BUF_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y82__R0_BUF_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R0_INV_0 (.A(tie_lo_T20Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y82__R1_BUF_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R1_INV_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R2_INV_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y82__R2_INV_1 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y82__R3_BUF_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y83__R0_BUF_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R0_INV_0 (.A(tie_lo_T20Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y83__R1_BUF_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R1_INV_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R2_INV_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y83__R2_INV_1 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y83__R3_BUF_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y84__R0_BUF_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R0_INV_0 (.A(tie_lo_T20Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y84__R1_BUF_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R1_INV_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R2_INV_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y84__R2_INV_1 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y84__R3_BUF_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y85__R0_BUF_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R0_INV_0 (.A(tie_lo_T20Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y85__R1_BUF_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R1_INV_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R2_INV_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y85__R2_INV_1 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y85__R3_BUF_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y86__R0_BUF_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R0_INV_0 (.A(tie_lo_T20Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y86__R1_BUF_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R1_INV_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R2_INV_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y86__R2_INV_1 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y86__R3_BUF_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y87__R0_BUF_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R0_INV_0 (.A(tie_lo_T20Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y87__R1_BUF_0 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R1_INV_0 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R2_INV_0 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y87__R2_INV_1 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y87__R3_BUF_0 (.A(tie_lo_T20Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y88__R0_BUF_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R0_INV_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y88__R1_BUF_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R1_INV_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R2_INV_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y88__R2_INV_1 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y88__R3_BUF_0 (.A(tie_lo_T20Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y89__R0_BUF_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R0_INV_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y89__R1_BUF_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R1_INV_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R2_INV_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y89__R2_INV_1 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y89__R3_BUF_0 (.A(tie_lo_T20Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y8__R0_BUF_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R0_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y8__R1_BUF_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R1_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R2_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y8__R2_INV_1 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y8__R3_BUF_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y9__R0_BUF_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R0_INV_0 (.A(tie_lo_T20Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y9__R1_BUF_0 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R1_INV_0 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T20Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R2_INV_0 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T20Y9__R2_INV_1 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T20Y9__R3_BUF_0 (.A(tie_lo_T20Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y0__R0_BUF_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R0_INV_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y0__R1_BUF_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R1_INV_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R2_INV_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y0__R2_INV_1 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y0__R3_BUF_0 (.A(tie_lo_T21Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y10__R0_BUF_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R0_INV_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y10__R1_BUF_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R1_INV_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R2_INV_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y10__R2_INV_1 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y10__R3_BUF_0 (.A(tie_lo_T21Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y11__R0_BUF_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R0_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y11__R1_BUF_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R1_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R2_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y11__R2_INV_1 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y11__R3_BUF_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y12__R0_BUF_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R0_INV_0 (.A(tie_lo_T21Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y12__R1_BUF_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R1_INV_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R2_INV_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y12__R2_INV_1 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y12__R3_BUF_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y13__R0_BUF_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R0_INV_0 (.A(tie_lo_T21Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y13__R1_BUF_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R1_INV_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R2_INV_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y13__R2_INV_1 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y13__R3_BUF_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y14__R0_BUF_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R0_INV_0 (.A(tie_lo_T21Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y14__R1_BUF_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R1_INV_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R2_INV_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y14__R2_INV_1 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y14__R3_BUF_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y15__R0_BUF_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R0_INV_0 (.A(tie_lo_T21Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y15__R1_BUF_0 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R1_INV_0 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R2_INV_0 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y15__R2_INV_1 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y15__R3_BUF_0 (.A(tie_lo_T21Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y16__R0_BUF_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R0_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y16__R1_BUF_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R1_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R2_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y16__R2_INV_1 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y16__R3_BUF_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y17__R0_BUF_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R0_INV_0 (.A(tie_lo_T21Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y17__R1_BUF_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R1_INV_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R2_INV_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y17__R2_INV_1 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y17__R3_BUF_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y18__R0_BUF_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R0_INV_0 (.A(tie_lo_T21Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y18__R1_BUF_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R1_INV_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R2_INV_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y18__R2_INV_1 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y18__R3_BUF_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y19__R0_BUF_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R0_INV_0 (.A(tie_lo_T21Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y19__R1_BUF_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R1_INV_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R2_INV_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y19__R2_INV_1 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y19__R3_BUF_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y1__R0_BUF_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R0_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y1__R1_BUF_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R1_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R2_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y1__R2_INV_1 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y1__R3_BUF_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y20__R0_BUF_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R0_INV_0 (.A(tie_lo_T21Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y20__R1_BUF_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R1_INV_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R2_INV_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y20__R2_INV_1 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y20__R3_BUF_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y21__R0_BUF_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R0_INV_0 (.A(tie_lo_T21Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y21__R1_BUF_0 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R1_INV_0 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R2_INV_0 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y21__R2_INV_1 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y21__R3_BUF_0 (.A(tie_lo_T21Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y22__R0_BUF_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R0_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y22__R1_BUF_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R1_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R2_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y22__R2_INV_1 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y22__R3_BUF_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y23__R0_BUF_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R0_INV_0 (.A(tie_lo_T21Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y23__R1_BUF_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R1_INV_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R2_INV_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y23__R2_INV_1 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y23__R3_BUF_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y24__R0_BUF_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R0_INV_0 (.A(tie_lo_T21Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y24__R1_BUF_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R1_INV_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R2_INV_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y24__R2_INV_1 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y24__R3_BUF_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y25__R0_BUF_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R0_INV_0 (.A(tie_lo_T21Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y25__R1_BUF_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R1_INV_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R2_INV_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y25__R2_INV_1 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y25__R3_BUF_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y26__R0_BUF_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R0_INV_0 (.A(tie_lo_T21Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y26__R1_BUF_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R1_INV_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R2_INV_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y26__R2_INV_1 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y26__R3_BUF_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y27__R0_BUF_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R0_INV_0 (.A(tie_lo_T21Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y27__R1_BUF_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R1_INV_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R2_INV_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y27__R2_INV_1 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y27__R3_BUF_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y28__R0_BUF_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R0_INV_0 (.A(tie_lo_T21Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y28__R1_BUF_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R1_INV_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R2_INV_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y28__R2_INV_1 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y28__R3_BUF_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y29__R0_BUF_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R0_INV_0 (.A(tie_lo_T21Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y29__R1_BUF_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R1_INV_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R2_INV_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y29__R2_INV_1 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y29__R3_BUF_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y2__R0_BUF_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R0_INV_0 (.A(tie_lo_T21Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y2__R1_BUF_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R1_INV_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R2_INV_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y2__R2_INV_1 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y2__R3_BUF_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y30__R0_BUF_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R0_INV_0 (.A(tie_lo_T21Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y30__R1_BUF_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R1_INV_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R2_INV_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y30__R2_INV_1 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y30__R3_BUF_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y31__R0_BUF_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R0_INV_0 (.A(tie_lo_T21Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y31__R1_BUF_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R1_INV_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R2_INV_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y31__R2_INV_1 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y31__R3_BUF_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y32__R0_BUF_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R0_INV_0 (.A(tie_lo_T21Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y32__R1_BUF_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R1_INV_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R2_INV_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y32__R2_INV_1 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y32__R3_BUF_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y33__R0_BUF_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R0_INV_0 (.A(tie_lo_T21Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y33__R1_BUF_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R1_INV_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R2_INV_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y33__R2_INV_1 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y33__R3_BUF_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y34__R0_BUF_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R0_INV_0 (.A(tie_lo_T21Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y34__R1_BUF_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R1_INV_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R2_INV_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y34__R2_INV_1 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y34__R3_BUF_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y35__R0_BUF_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R0_INV_0 (.A(tie_lo_T21Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y35__R1_BUF_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R1_INV_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R2_INV_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y35__R2_INV_1 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y35__R3_BUF_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y36__R0_BUF_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R0_INV_0 (.A(tie_lo_T21Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y36__R1_BUF_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R1_INV_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R2_INV_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y36__R2_INV_1 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y36__R3_BUF_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y37__R0_BUF_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R0_INV_0 (.A(tie_lo_T21Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y37__R1_BUF_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R1_INV_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R2_INV_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y37__R2_INV_1 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y37__R3_BUF_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y38__R0_BUF_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R0_INV_0 (.A(tie_lo_T21Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y38__R1_BUF_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R1_INV_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R2_INV_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y38__R2_INV_1 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y38__R3_BUF_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y39__R0_BUF_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R0_INV_0 (.A(tie_lo_T21Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y39__R1_BUF_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R1_INV_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R2_INV_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y39__R2_INV_1 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y39__R3_BUF_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y3__R0_BUF_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R0_INV_0 (.A(tie_lo_T21Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y3__R1_BUF_0 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R1_INV_0 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R2_INV_0 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y3__R2_INV_1 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y3__R3_BUF_0 (.A(tie_lo_T21Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y40__R0_BUF_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R0_INV_0 (.A(tie_lo_T21Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y40__R1_BUF_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R1_INV_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R2_INV_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y40__R2_INV_1 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y40__R3_BUF_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y41__R0_BUF_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R0_INV_0 (.A(tie_lo_T21Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y41__R1_BUF_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R1_INV_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R2_INV_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y41__R2_INV_1 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y41__R3_BUF_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y42__R0_BUF_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R0_INV_0 (.A(tie_lo_T21Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y42__R1_BUF_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R1_INV_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R2_INV_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y42__R2_INV_1 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y42__R3_BUF_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y43__R0_BUF_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R0_INV_0 (.A(tie_lo_T21Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y43__R1_BUF_0 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R1_INV_0 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R2_INV_0 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y43__R2_INV_1 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y43__R3_BUF_0 (.A(tie_lo_T21Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y44__R0_BUF_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R0_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y44__R1_BUF_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R1_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R2_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y44__R2_INV_1 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y44__R3_BUF_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y45__R0_BUF_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R0_INV_0 (.A(tie_lo_T21Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y45__R1_BUF_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R1_INV_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R2_INV_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y45__R2_INV_1 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y45__R3_BUF_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y46__R0_BUF_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R0_INV_0 (.A(tie_lo_T21Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y46__R1_BUF_0 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R1_INV_0 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R2_INV_0 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y46__R2_INV_1 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y46__R3_BUF_0 (.A(tie_lo_T21Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y47__R0_BUF_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R0_INV_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y47__R1_BUF_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R1_INV_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R2_INV_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y47__R2_INV_1 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y47__R3_BUF_0 (.A(tie_lo_T21Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y48__R0_BUF_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R0_INV_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y48__R1_BUF_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R1_INV_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R2_INV_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y48__R2_INV_1 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y48__R3_BUF_0 (.A(tie_lo_T21Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y49__R0_BUF_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R0_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y49__R1_BUF_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R1_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R2_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y49__R2_INV_1 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y49__R3_BUF_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y4__R0_BUF_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R0_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y4__R1_BUF_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R1_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R2_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y4__R2_INV_1 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y4__R3_BUF_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y50__R0_BUF_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R0_INV_0 (.A(tie_lo_T21Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y50__R1_BUF_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R1_INV_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R2_INV_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y50__R2_INV_1 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y50__R3_BUF_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y51__R0_BUF_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R0_INV_0 (.A(tie_lo_T21Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y51__R1_BUF_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R1_INV_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R2_INV_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y51__R2_INV_1 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y51__R3_BUF_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y52__R0_BUF_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R0_INV_0 (.A(tie_lo_T21Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y52__R1_BUF_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R1_INV_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R2_INV_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y52__R2_INV_1 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y52__R3_BUF_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y53__R0_BUF_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R0_INV_0 (.A(tie_lo_T21Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y53__R1_BUF_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R1_INV_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R2_INV_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y53__R2_INV_1 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y53__R3_BUF_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y54__R0_BUF_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R0_INV_0 (.A(tie_lo_T21Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y54__R1_BUF_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R1_INV_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R2_INV_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y54__R2_INV_1 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y54__R3_BUF_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y55__R0_BUF_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R0_INV_0 (.A(tie_lo_T21Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y55__R1_BUF_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R1_INV_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R2_INV_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y55__R2_INV_1 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y55__R3_BUF_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y56__R0_BUF_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R0_INV_0 (.A(tie_lo_T21Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y56__R1_BUF_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R1_INV_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R2_INV_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y56__R2_INV_1 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y56__R3_BUF_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y57__R0_BUF_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R0_INV_0 (.A(tie_lo_T21Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y57__R1_BUF_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R1_INV_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R2_INV_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y57__R2_INV_1 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y57__R3_BUF_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y58__R0_BUF_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R0_INV_0 (.A(tie_lo_T21Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y58__R1_BUF_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R1_INV_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R2_INV_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y58__R2_INV_1 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y58__R3_BUF_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y59__R0_BUF_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R0_INV_0 (.A(tie_lo_T21Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y59__R1_BUF_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R1_INV_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R2_INV_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y59__R2_INV_1 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y59__R3_BUF_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y5__R0_BUF_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R0_INV_0 (.A(tie_lo_T21Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y5__R1_BUF_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R1_INV_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R2_INV_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y5__R2_INV_1 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y5__R3_BUF_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y60__R0_BUF_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R0_INV_0 (.A(tie_lo_T21Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y60__R1_BUF_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R1_INV_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R2_INV_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y60__R2_INV_1 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y60__R3_BUF_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y61__R0_BUF_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R0_INV_0 (.A(tie_lo_T21Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y61__R1_BUF_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R1_INV_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R2_INV_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y61__R2_INV_1 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y61__R3_BUF_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y62__R0_BUF_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R0_INV_0 (.A(tie_lo_T21Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y62__R1_BUF_0 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R1_INV_0 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R2_INV_0 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y62__R2_INV_1 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y62__R3_BUF_0 (.A(tie_lo_T21Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y63__R0_BUF_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R0_INV_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y63__R1_BUF_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R1_INV_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R2_INV_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y63__R2_INV_1 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y63__R3_BUF_0 (.A(tie_lo_T21Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y64__R0_BUF_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R0_INV_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y64__R1_BUF_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R1_INV_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R2_INV_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y64__R2_INV_1 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y64__R3_BUF_0 (.A(tie_lo_T21Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y65__R0_BUF_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R0_INV_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y65__R1_BUF_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R1_INV_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R2_INV_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y65__R2_INV_1 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y65__R3_BUF_0 (.A(tie_lo_T21Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y66__R0_BUF_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R0_INV_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y66__R1_BUF_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R1_INV_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R2_INV_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y66__R2_INV_1 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y66__R3_BUF_0 (.A(tie_lo_T21Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y67__R0_BUF_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R0_INV_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y67__R1_BUF_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R1_INV_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R2_INV_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y67__R2_INV_1 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y67__R3_BUF_0 (.A(tie_lo_T21Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y68__R0_BUF_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R0_INV_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y68__R1_BUF_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R1_INV_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R2_INV_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y68__R2_INV_1 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y68__R3_BUF_0 (.A(tie_lo_T21Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y69__R0_BUF_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R0_INV_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y69__R1_BUF_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R1_INV_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R2_INV_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y69__R2_INV_1 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y69__R3_BUF_0 (.A(tie_lo_T21Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y6__R0_BUF_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R0_INV_0 (.A(tie_lo_T21Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y6__R1_BUF_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R1_INV_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R2_INV_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y6__R2_INV_1 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y6__R3_BUF_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y70__R0_BUF_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R0_INV_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y70__R1_BUF_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R1_INV_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R2_INV_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y70__R2_INV_1 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y70__R3_BUF_0 (.A(tie_lo_T21Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y71__R0_BUF_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R0_INV_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y71__R1_BUF_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R1_INV_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R2_INV_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y71__R2_INV_1 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y71__R3_BUF_0 (.A(tie_lo_T21Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y72__R0_BUF_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R0_INV_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y72__R1_BUF_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R1_INV_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R2_INV_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y72__R2_INV_1 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y72__R3_BUF_0 (.A(tie_lo_T21Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y73__R0_BUF_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R0_INV_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y73__R1_BUF_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R1_INV_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R2_INV_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y73__R2_INV_1 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y73__R3_BUF_0 (.A(tie_lo_T21Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y74__R0_BUF_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R0_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y74__R1_BUF_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R1_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R2_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y74__R2_INV_1 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y74__R3_BUF_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y75__R0_BUF_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R0_INV_0 (.A(tie_lo_T21Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y75__R1_BUF_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R1_INV_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R2_INV_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y75__R2_INV_1 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y75__R3_BUF_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y76__R0_BUF_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R0_INV_0 (.A(tie_lo_T21Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y76__R1_BUF_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R1_INV_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R2_INV_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y76__R2_INV_1 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y76__R3_BUF_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y77__R0_BUF_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R0_INV_0 (.A(tie_lo_T21Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y77__R1_BUF_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R1_INV_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R2_INV_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y77__R2_INV_1 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y77__R3_BUF_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y78__R0_BUF_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R0_INV_0 (.A(tie_lo_T21Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y78__R1_BUF_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R1_INV_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R2_INV_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y78__R2_INV_1 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y78__R3_BUF_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y79__R0_BUF_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R0_INV_0 (.A(tie_lo_T21Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y79__R1_BUF_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R1_INV_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R2_INV_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y79__R2_INV_1 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y79__R3_BUF_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y7__R0_BUF_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R0_INV_0 (.A(tie_lo_T21Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y7__R1_BUF_0 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R1_INV_0 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R2_INV_0 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y7__R2_INV_1 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y7__R3_BUF_0 (.A(tie_lo_T21Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y80__R0_BUF_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R0_INV_0 (.A(tie_lo_T21Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y80__R1_BUF_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R1_INV_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R2_INV_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y80__R2_INV_1 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y80__R3_BUF_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y81__R0_BUF_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R0_INV_0 (.A(tie_lo_T21Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y81__R1_BUF_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R1_INV_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R2_INV_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y81__R2_INV_1 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y81__R3_BUF_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y82__R0_BUF_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R0_INV_0 (.A(tie_lo_T21Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y82__R1_BUF_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R1_INV_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R2_INV_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y82__R2_INV_1 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y82__R3_BUF_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y83__R0_BUF_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R0_INV_0 (.A(tie_lo_T21Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y83__R1_BUF_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R1_INV_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R2_INV_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y83__R2_INV_1 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y83__R3_BUF_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y84__R0_BUF_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R0_INV_0 (.A(tie_lo_T21Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y84__R1_BUF_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R1_INV_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R2_INV_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y84__R2_INV_1 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y84__R3_BUF_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y85__R0_BUF_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R0_INV_0 (.A(tie_lo_T21Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y85__R1_BUF_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R1_INV_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R2_INV_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y85__R2_INV_1 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y85__R3_BUF_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y86__R0_BUF_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R0_INV_0 (.A(tie_lo_T21Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y86__R1_BUF_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R1_INV_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R2_INV_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y86__R2_INV_1 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y86__R3_BUF_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y87__R0_BUF_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R0_INV_0 (.A(tie_lo_T21Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y87__R1_BUF_0 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R1_INV_0 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R2_INV_0 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y87__R2_INV_1 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y87__R3_BUF_0 (.A(tie_lo_T21Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y88__R0_BUF_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R0_INV_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y88__R1_BUF_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R1_INV_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R2_INV_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y88__R2_INV_1 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y88__R3_BUF_0 (.A(tie_lo_T21Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y89__R0_BUF_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R0_INV_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y89__R1_BUF_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R1_INV_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R2_INV_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y89__R2_INV_1 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y89__R3_BUF_0 (.A(tie_lo_T21Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y8__R0_BUF_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R0_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y8__R1_BUF_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R1_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R2_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y8__R2_INV_1 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y8__R3_BUF_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y9__R0_BUF_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R0_INV_0 (.A(tie_lo_T21Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y9__R1_BUF_0 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R1_INV_0 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T21Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R2_INV_0 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T21Y9__R2_INV_1 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T21Y9__R3_BUF_0 (.A(tie_lo_T21Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y0__R0_BUF_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R0_INV_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y0__R1_BUF_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R1_INV_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R2_INV_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y0__R2_INV_1 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y0__R3_BUF_0 (.A(tie_lo_T22Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y10__R0_BUF_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R0_INV_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y10__R1_BUF_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R1_INV_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R2_INV_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y10__R2_INV_1 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y10__R3_BUF_0 (.A(tie_lo_T22Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y11__R0_BUF_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R0_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y11__R1_BUF_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R1_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R2_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y11__R2_INV_1 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y11__R3_BUF_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y12__R0_BUF_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R0_INV_0 (.A(tie_lo_T22Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y12__R1_BUF_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R1_INV_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R2_INV_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y12__R2_INV_1 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y12__R3_BUF_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y13__R0_BUF_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R0_INV_0 (.A(tie_lo_T22Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y13__R1_BUF_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R1_INV_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R2_INV_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y13__R2_INV_1 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y13__R3_BUF_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y14__R0_BUF_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R0_INV_0 (.A(tie_lo_T22Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y14__R1_BUF_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R1_INV_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R2_INV_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y14__R2_INV_1 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y14__R3_BUF_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y15__R0_BUF_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R0_INV_0 (.A(tie_lo_T22Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y15__R1_BUF_0 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R1_INV_0 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R2_INV_0 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y15__R2_INV_1 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y15__R3_BUF_0 (.A(tie_lo_T22Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y16__R0_BUF_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R0_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y16__R1_BUF_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R1_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R2_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y16__R2_INV_1 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y16__R3_BUF_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y17__R0_BUF_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R0_INV_0 (.A(tie_lo_T22Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y17__R1_BUF_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R1_INV_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R2_INV_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y17__R2_INV_1 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y17__R3_BUF_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y18__R0_BUF_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R0_INV_0 (.A(tie_lo_T22Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y18__R1_BUF_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R1_INV_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R2_INV_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y18__R2_INV_1 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y18__R3_BUF_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y19__R0_BUF_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R0_INV_0 (.A(tie_lo_T22Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y19__R1_BUF_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R1_INV_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R2_INV_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y19__R2_INV_1 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y19__R3_BUF_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y1__R0_BUF_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R0_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y1__R1_BUF_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R1_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R2_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y1__R2_INV_1 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y1__R3_BUF_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y20__R0_BUF_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R0_INV_0 (.A(tie_lo_T22Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y20__R1_BUF_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R1_INV_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R2_INV_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y20__R2_INV_1 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y20__R3_BUF_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y21__R0_BUF_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R0_INV_0 (.A(tie_lo_T22Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y21__R1_BUF_0 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R1_INV_0 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R2_INV_0 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y21__R2_INV_1 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y21__R3_BUF_0 (.A(tie_lo_T22Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y22__R0_BUF_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R0_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y22__R1_BUF_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R1_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R2_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y22__R2_INV_1 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y22__R3_BUF_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y23__R0_BUF_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R0_INV_0 (.A(tie_lo_T22Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y23__R1_BUF_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R1_INV_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R2_INV_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y23__R2_INV_1 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y23__R3_BUF_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y24__R0_BUF_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R0_INV_0 (.A(tie_lo_T22Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y24__R1_BUF_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R1_INV_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R2_INV_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y24__R2_INV_1 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y24__R3_BUF_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y25__R0_BUF_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R0_INV_0 (.A(tie_lo_T22Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y25__R1_BUF_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R1_INV_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R2_INV_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y25__R2_INV_1 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y25__R3_BUF_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y26__R0_BUF_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R0_INV_0 (.A(tie_lo_T22Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y26__R1_BUF_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R1_INV_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R2_INV_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y26__R2_INV_1 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y26__R3_BUF_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y27__R0_BUF_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R0_INV_0 (.A(tie_lo_T22Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y27__R1_BUF_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R1_INV_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R2_INV_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y27__R2_INV_1 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y27__R3_BUF_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y28__R0_BUF_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R0_INV_0 (.A(tie_lo_T22Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y28__R1_BUF_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R1_INV_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R2_INV_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y28__R2_INV_1 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y28__R3_BUF_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y29__R0_BUF_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R0_INV_0 (.A(tie_lo_T22Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y29__R1_BUF_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R1_INV_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R2_INV_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y29__R2_INV_1 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y29__R3_BUF_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y2__R0_BUF_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R0_INV_0 (.A(tie_lo_T22Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y2__R1_BUF_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R1_INV_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R2_INV_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y2__R2_INV_1 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y2__R3_BUF_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y30__R0_BUF_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R0_INV_0 (.A(tie_lo_T22Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y30__R1_BUF_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R1_INV_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R2_INV_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y30__R2_INV_1 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y30__R3_BUF_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y31__R0_BUF_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R0_INV_0 (.A(tie_lo_T22Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y31__R1_BUF_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R1_INV_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R2_INV_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y31__R2_INV_1 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y31__R3_BUF_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y32__R0_BUF_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R0_INV_0 (.A(tie_lo_T22Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y32__R1_BUF_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R1_INV_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R2_INV_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y32__R2_INV_1 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y32__R3_BUF_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y33__R0_BUF_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R0_INV_0 (.A(tie_lo_T22Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y33__R1_BUF_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R1_INV_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R2_INV_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y33__R2_INV_1 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y33__R3_BUF_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y34__R0_BUF_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R0_INV_0 (.A(tie_lo_T22Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y34__R1_BUF_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R1_INV_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R2_INV_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y34__R2_INV_1 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y34__R3_BUF_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y35__R0_BUF_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R0_INV_0 (.A(tie_lo_T22Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y35__R1_BUF_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R1_INV_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R2_INV_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y35__R2_INV_1 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y35__R3_BUF_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y36__R0_BUF_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R0_INV_0 (.A(tie_lo_T22Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y36__R1_BUF_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R1_INV_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R2_INV_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y36__R2_INV_1 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y36__R3_BUF_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y37__R0_BUF_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R0_INV_0 (.A(tie_lo_T22Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y37__R1_BUF_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R1_INV_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R2_INV_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y37__R2_INV_1 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y37__R3_BUF_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y38__R0_BUF_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R0_INV_0 (.A(tie_lo_T22Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y38__R1_BUF_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R1_INV_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R2_INV_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y38__R2_INV_1 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y38__R3_BUF_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y39__R0_BUF_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R0_INV_0 (.A(tie_lo_T22Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y39__R1_BUF_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R1_INV_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R2_INV_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y39__R2_INV_1 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y39__R3_BUF_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y3__R0_BUF_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R0_INV_0 (.A(tie_lo_T22Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y3__R1_BUF_0 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R1_INV_0 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R2_INV_0 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y3__R2_INV_1 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y3__R3_BUF_0 (.A(tie_lo_T22Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y40__R0_BUF_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R0_INV_0 (.A(tie_lo_T22Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y40__R1_BUF_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R1_INV_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R2_INV_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y40__R2_INV_1 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y40__R3_BUF_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y41__R0_BUF_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R0_INV_0 (.A(tie_lo_T22Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y41__R1_BUF_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R1_INV_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R2_INV_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y41__R2_INV_1 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y41__R3_BUF_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y42__R0_BUF_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R0_INV_0 (.A(tie_lo_T22Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y42__R1_BUF_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R1_INV_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R2_INV_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y42__R2_INV_1 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y42__R3_BUF_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y43__R0_BUF_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R0_INV_0 (.A(tie_lo_T22Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y43__R1_BUF_0 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R1_INV_0 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R2_INV_0 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y43__R2_INV_1 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y43__R3_BUF_0 (.A(tie_lo_T22Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y44__R0_BUF_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R0_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y44__R1_BUF_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R1_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R2_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y44__R2_INV_1 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y44__R3_BUF_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y45__R0_BUF_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R0_INV_0 (.A(tie_lo_T22Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y45__R1_BUF_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R1_INV_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R2_INV_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y45__R2_INV_1 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y45__R3_BUF_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y46__R0_BUF_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R0_INV_0 (.A(tie_lo_T22Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y46__R1_BUF_0 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R1_INV_0 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R2_INV_0 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y46__R2_INV_1 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y46__R3_BUF_0 (.A(tie_lo_T22Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y47__R0_BUF_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R0_INV_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y47__R1_BUF_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R1_INV_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R2_INV_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y47__R2_INV_1 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y47__R3_BUF_0 (.A(tie_lo_T22Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y48__R0_BUF_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R0_INV_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y48__R1_BUF_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R1_INV_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R2_INV_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y48__R2_INV_1 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y48__R3_BUF_0 (.A(tie_lo_T22Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y49__R0_BUF_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R0_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y49__R1_BUF_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R1_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R2_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y49__R2_INV_1 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y49__R3_BUF_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y4__R0_BUF_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R0_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y4__R1_BUF_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R1_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R2_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y4__R2_INV_1 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y4__R3_BUF_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y50__R0_BUF_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R0_INV_0 (.A(tie_lo_T22Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y50__R1_BUF_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R1_INV_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R2_INV_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y50__R2_INV_1 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y50__R3_BUF_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y51__R0_BUF_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R0_INV_0 (.A(tie_lo_T22Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y51__R1_BUF_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R1_INV_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R2_INV_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y51__R2_INV_1 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y51__R3_BUF_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y52__R0_BUF_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R0_INV_0 (.A(tie_lo_T22Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y52__R1_BUF_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R1_INV_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R2_INV_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y52__R2_INV_1 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y52__R3_BUF_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y53__R0_BUF_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R0_INV_0 (.A(tie_lo_T22Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y53__R1_BUF_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R1_INV_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R2_INV_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y53__R2_INV_1 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y53__R3_BUF_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y54__R0_BUF_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R0_INV_0 (.A(tie_lo_T22Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y54__R1_BUF_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R1_INV_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R2_INV_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y54__R2_INV_1 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y54__R3_BUF_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y55__R0_BUF_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R0_INV_0 (.A(tie_lo_T22Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y55__R1_BUF_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R1_INV_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R2_INV_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y55__R2_INV_1 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y55__R3_BUF_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y56__R0_BUF_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R0_INV_0 (.A(tie_lo_T22Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y56__R1_BUF_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R1_INV_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R2_INV_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y56__R2_INV_1 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y56__R3_BUF_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y57__R0_BUF_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R0_INV_0 (.A(tie_lo_T22Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y57__R1_BUF_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R1_INV_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R2_INV_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y57__R2_INV_1 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y57__R3_BUF_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y58__R0_BUF_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R0_INV_0 (.A(tie_lo_T22Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y58__R1_BUF_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R1_INV_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R2_INV_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y58__R2_INV_1 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y58__R3_BUF_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y59__R0_BUF_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R0_INV_0 (.A(tie_lo_T22Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y59__R1_BUF_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R1_INV_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R2_INV_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y59__R2_INV_1 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y59__R3_BUF_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y5__R0_BUF_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R0_INV_0 (.A(tie_lo_T22Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y5__R1_BUF_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R1_INV_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R2_INV_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y5__R2_INV_1 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y5__R3_BUF_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y60__R0_BUF_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R0_INV_0 (.A(tie_lo_T22Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y60__R1_BUF_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R1_INV_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R2_INV_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y60__R2_INV_1 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y60__R3_BUF_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y61__R0_BUF_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R0_INV_0 (.A(tie_lo_T22Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y61__R1_BUF_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R1_INV_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R2_INV_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y61__R2_INV_1 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y61__R3_BUF_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y62__R0_BUF_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R0_INV_0 (.A(tie_lo_T22Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y62__R1_BUF_0 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R1_INV_0 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R2_INV_0 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y62__R2_INV_1 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y62__R3_BUF_0 (.A(tie_lo_T22Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y63__R0_BUF_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R0_INV_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y63__R1_BUF_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R1_INV_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R2_INV_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y63__R2_INV_1 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y63__R3_BUF_0 (.A(tie_lo_T22Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y64__R0_BUF_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R0_INV_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y64__R1_BUF_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R1_INV_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R2_INV_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y64__R2_INV_1 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y64__R3_BUF_0 (.A(tie_lo_T22Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y65__R0_BUF_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R0_INV_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y65__R1_BUF_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R1_INV_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R2_INV_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y65__R2_INV_1 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y65__R3_BUF_0 (.A(tie_lo_T22Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y66__R0_BUF_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R0_INV_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y66__R1_BUF_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R1_INV_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R2_INV_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y66__R2_INV_1 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y66__R3_BUF_0 (.A(tie_lo_T22Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y67__R0_BUF_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R0_INV_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y67__R1_BUF_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R1_INV_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R2_INV_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y67__R2_INV_1 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y67__R3_BUF_0 (.A(tie_lo_T22Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y68__R0_BUF_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R0_INV_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y68__R1_BUF_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R1_INV_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R2_INV_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y68__R2_INV_1 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y68__R3_BUF_0 (.A(tie_lo_T22Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y69__R0_BUF_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R0_INV_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y69__R1_BUF_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R1_INV_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R2_INV_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y69__R2_INV_1 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y69__R3_BUF_0 (.A(tie_lo_T22Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y6__R0_BUF_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R0_INV_0 (.A(tie_lo_T22Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y6__R1_BUF_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R1_INV_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R2_INV_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y6__R2_INV_1 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y6__R3_BUF_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y70__R0_BUF_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R0_INV_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y70__R1_BUF_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R1_INV_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R2_INV_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y70__R2_INV_1 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y70__R3_BUF_0 (.A(tie_lo_T22Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y71__R0_BUF_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R0_INV_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y71__R1_BUF_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R1_INV_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R2_INV_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y71__R2_INV_1 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y71__R3_BUF_0 (.A(tie_lo_T22Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y72__R0_BUF_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R0_INV_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y72__R1_BUF_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R1_INV_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R2_INV_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y72__R2_INV_1 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y72__R3_BUF_0 (.A(tie_lo_T22Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y73__R0_BUF_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R0_INV_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y73__R1_BUF_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R1_INV_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R2_INV_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y73__R2_INV_1 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y73__R3_BUF_0 (.A(tie_lo_T22Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y74__R0_BUF_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R0_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y74__R1_BUF_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R1_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R2_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y74__R2_INV_1 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y74__R3_BUF_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y75__R0_BUF_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R0_INV_0 (.A(tie_lo_T22Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y75__R1_BUF_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R1_INV_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R2_INV_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y75__R2_INV_1 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y75__R3_BUF_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y76__R0_BUF_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R0_INV_0 (.A(tie_lo_T22Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y76__R1_BUF_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R1_INV_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R2_INV_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y76__R2_INV_1 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y76__R3_BUF_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y77__R0_BUF_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R0_INV_0 (.A(tie_lo_T22Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y77__R1_BUF_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R1_INV_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R2_INV_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y77__R2_INV_1 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y77__R3_BUF_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y78__R0_BUF_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R0_INV_0 (.A(tie_lo_T22Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y78__R1_BUF_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R1_INV_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R2_INV_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y78__R2_INV_1 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y78__R3_BUF_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y79__R0_BUF_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R0_INV_0 (.A(tie_lo_T22Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y79__R1_BUF_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R1_INV_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R2_INV_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y79__R2_INV_1 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y79__R3_BUF_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y7__R0_BUF_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R0_INV_0 (.A(tie_lo_T22Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y7__R1_BUF_0 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R1_INV_0 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R2_INV_0 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y7__R2_INV_1 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y7__R3_BUF_0 (.A(tie_lo_T22Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y80__R0_BUF_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R0_INV_0 (.A(tie_lo_T22Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y80__R1_BUF_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R1_INV_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R2_INV_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y80__R2_INV_1 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y80__R3_BUF_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y81__R0_BUF_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R0_INV_0 (.A(tie_lo_T22Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y81__R1_BUF_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R1_INV_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R2_INV_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y81__R2_INV_1 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y81__R3_BUF_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y82__R0_BUF_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R0_INV_0 (.A(tie_lo_T22Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y82__R1_BUF_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R1_INV_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R2_INV_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y82__R2_INV_1 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y82__R3_BUF_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y83__R0_BUF_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R0_INV_0 (.A(tie_lo_T22Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y83__R1_BUF_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R1_INV_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R2_INV_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y83__R2_INV_1 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y83__R3_BUF_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y84__R0_BUF_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R0_INV_0 (.A(tie_lo_T22Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y84__R1_BUF_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R1_INV_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R2_INV_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y84__R2_INV_1 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y84__R3_BUF_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y85__R0_BUF_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R0_INV_0 (.A(tie_lo_T22Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y85__R1_BUF_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R1_INV_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R2_INV_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y85__R2_INV_1 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y85__R3_BUF_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y86__R0_BUF_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R0_INV_0 (.A(tie_lo_T22Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y86__R1_BUF_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R1_INV_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R2_INV_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y86__R2_INV_1 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y86__R3_BUF_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y87__R0_BUF_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R0_INV_0 (.A(tie_lo_T22Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y87__R1_BUF_0 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R1_INV_0 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R2_INV_0 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y87__R2_INV_1 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y87__R3_BUF_0 (.A(tie_lo_T22Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y88__R0_BUF_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R0_INV_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y88__R1_BUF_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R1_INV_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R2_INV_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y88__R2_INV_1 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y88__R3_BUF_0 (.A(tie_lo_T22Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y89__R0_BUF_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R0_INV_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y89__R1_BUF_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R1_INV_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R2_INV_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y89__R2_INV_1 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y89__R3_BUF_0 (.A(tie_lo_T22Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y8__R0_BUF_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R0_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y8__R1_BUF_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R1_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R2_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y8__R2_INV_1 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y8__R3_BUF_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y9__R0_BUF_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R0_INV_0 (.A(tie_lo_T22Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y9__R1_BUF_0 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R1_INV_0 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T22Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R2_INV_0 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T22Y9__R2_INV_1 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T22Y9__R3_BUF_0 (.A(tie_lo_T22Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y0__R0_BUF_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R0_INV_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y0__R1_BUF_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R1_INV_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R2_INV_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y0__R2_INV_1 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y0__R3_BUF_0 (.A(tie_lo_T23Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y10__R0_BUF_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R0_INV_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y10__R1_BUF_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R1_INV_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R2_INV_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y10__R2_INV_1 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y10__R3_BUF_0 (.A(tie_lo_T23Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y11__R0_BUF_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R0_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y11__R1_BUF_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R1_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R2_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y11__R2_INV_1 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y11__R3_BUF_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y12__R0_BUF_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R0_INV_0 (.A(tie_lo_T23Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y12__R1_BUF_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R1_INV_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R2_INV_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y12__R2_INV_1 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y12__R3_BUF_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y13__R0_BUF_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R0_INV_0 (.A(tie_lo_T23Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y13__R1_BUF_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R1_INV_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R2_INV_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y13__R2_INV_1 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y13__R3_BUF_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y14__R0_BUF_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R0_INV_0 (.A(tie_lo_T23Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y14__R1_BUF_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R1_INV_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R2_INV_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y14__R2_INV_1 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y14__R3_BUF_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y15__R0_BUF_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R0_INV_0 (.A(tie_lo_T23Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y15__R1_BUF_0 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R1_INV_0 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R2_INV_0 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y15__R2_INV_1 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y15__R3_BUF_0 (.A(tie_lo_T23Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y16__R0_BUF_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R0_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y16__R1_BUF_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R1_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R2_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y16__R2_INV_1 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y16__R3_BUF_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y17__R0_BUF_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R0_INV_0 (.A(tie_lo_T23Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y17__R1_BUF_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R1_INV_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R2_INV_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y17__R2_INV_1 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y17__R3_BUF_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y18__R0_BUF_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R0_INV_0 (.A(tie_lo_T23Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y18__R1_BUF_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R1_INV_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R2_INV_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y18__R2_INV_1 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y18__R3_BUF_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y19__R0_BUF_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R0_INV_0 (.A(tie_lo_T23Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y19__R1_BUF_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R1_INV_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R2_INV_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y19__R2_INV_1 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y19__R3_BUF_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y1__R0_BUF_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R0_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y1__R1_BUF_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R1_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R2_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y1__R2_INV_1 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y1__R3_BUF_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y20__R0_BUF_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R0_INV_0 (.A(tie_lo_T23Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y20__R1_BUF_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R1_INV_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R2_INV_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y20__R2_INV_1 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y20__R3_BUF_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y21__R0_BUF_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R0_INV_0 (.A(tie_lo_T23Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y21__R1_BUF_0 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R1_INV_0 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R2_INV_0 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y21__R2_INV_1 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y21__R3_BUF_0 (.A(tie_lo_T23Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y22__R0_BUF_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R0_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y22__R1_BUF_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R1_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R2_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y22__R2_INV_1 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y22__R3_BUF_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y23__R0_BUF_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R0_INV_0 (.A(tie_lo_T23Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y23__R1_BUF_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R1_INV_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R2_INV_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y23__R2_INV_1 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y23__R3_BUF_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y24__R0_BUF_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R0_INV_0 (.A(tie_lo_T23Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y24__R1_BUF_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R1_INV_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R2_INV_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y24__R2_INV_1 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y24__R3_BUF_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y25__R0_BUF_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R0_INV_0 (.A(tie_lo_T23Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y25__R1_BUF_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R1_INV_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R2_INV_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y25__R2_INV_1 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y25__R3_BUF_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y26__R0_BUF_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R0_INV_0 (.A(tie_lo_T23Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y26__R1_BUF_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R1_INV_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R2_INV_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y26__R2_INV_1 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y26__R3_BUF_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y27__R0_BUF_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R0_INV_0 (.A(tie_lo_T23Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y27__R1_BUF_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R1_INV_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R2_INV_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y27__R2_INV_1 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y27__R3_BUF_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y28__R0_BUF_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R0_INV_0 (.A(tie_lo_T23Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y28__R1_BUF_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R1_INV_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R2_INV_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y28__R2_INV_1 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y28__R3_BUF_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y29__R0_BUF_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R0_INV_0 (.A(tie_lo_T23Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y29__R1_BUF_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R1_INV_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R2_INV_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y29__R2_INV_1 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y29__R3_BUF_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y2__R0_BUF_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R0_INV_0 (.A(tie_lo_T23Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y2__R1_BUF_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R1_INV_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R2_INV_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y2__R2_INV_1 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y2__R3_BUF_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y30__R0_BUF_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R0_INV_0 (.A(tie_lo_T23Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y30__R1_BUF_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R1_INV_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R2_INV_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y30__R2_INV_1 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y30__R3_BUF_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y31__R0_BUF_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R0_INV_0 (.A(tie_lo_T23Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y31__R1_BUF_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R1_INV_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R2_INV_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y31__R2_INV_1 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y31__R3_BUF_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y32__R0_BUF_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R0_INV_0 (.A(tie_lo_T23Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y32__R1_BUF_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R1_INV_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R2_INV_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y32__R2_INV_1 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y32__R3_BUF_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y33__R0_BUF_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R0_INV_0 (.A(tie_lo_T23Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y33__R1_BUF_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R1_INV_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R2_INV_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y33__R2_INV_1 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y33__R3_BUF_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y34__R0_BUF_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R0_INV_0 (.A(tie_lo_T23Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y34__R1_BUF_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R1_INV_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R2_INV_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y34__R2_INV_1 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y34__R3_BUF_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y35__R0_BUF_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R0_INV_0 (.A(tie_lo_T23Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y35__R1_BUF_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R1_INV_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R2_INV_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y35__R2_INV_1 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y35__R3_BUF_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y36__R0_BUF_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R0_INV_0 (.A(tie_lo_T23Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y36__R1_BUF_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R1_INV_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R2_INV_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y36__R2_INV_1 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y36__R3_BUF_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y37__R0_BUF_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R0_INV_0 (.A(tie_lo_T23Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y37__R1_BUF_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R1_INV_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R2_INV_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y37__R2_INV_1 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y37__R3_BUF_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y38__R0_BUF_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R0_INV_0 (.A(tie_lo_T23Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y38__R1_BUF_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R1_INV_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R2_INV_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y38__R2_INV_1 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y38__R3_BUF_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y39__R0_BUF_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R0_INV_0 (.A(tie_lo_T23Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y39__R1_BUF_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R1_INV_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R2_INV_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y39__R2_INV_1 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y39__R3_BUF_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y3__R0_BUF_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R0_INV_0 (.A(tie_lo_T23Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y3__R1_BUF_0 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R1_INV_0 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R2_INV_0 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y3__R2_INV_1 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y3__R3_BUF_0 (.A(tie_lo_T23Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y40__R0_BUF_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R0_INV_0 (.A(tie_lo_T23Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y40__R1_BUF_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R1_INV_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R2_INV_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y40__R2_INV_1 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y40__R3_BUF_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y41__R0_BUF_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R0_INV_0 (.A(tie_lo_T23Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y41__R1_BUF_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R1_INV_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R2_INV_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y41__R2_INV_1 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y41__R3_BUF_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y42__R0_BUF_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R0_INV_0 (.A(tie_lo_T23Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y42__R1_BUF_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R1_INV_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R2_INV_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y42__R2_INV_1 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y42__R3_BUF_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y43__R0_BUF_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R0_INV_0 (.A(tie_lo_T23Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y43__R1_BUF_0 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R1_INV_0 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R2_INV_0 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y43__R2_INV_1 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y43__R3_BUF_0 (.A(tie_lo_T23Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y44__R0_BUF_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R0_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y44__R1_BUF_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R1_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R2_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y44__R2_INV_1 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y44__R3_BUF_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y45__R0_BUF_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R0_INV_0 (.A(tie_lo_T23Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y45__R1_BUF_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R1_INV_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R2_INV_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y45__R2_INV_1 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y45__R3_BUF_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y46__R0_BUF_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R0_INV_0 (.A(tie_lo_T23Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y46__R1_BUF_0 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R1_INV_0 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R2_INV_0 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y46__R2_INV_1 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y46__R3_BUF_0 (.A(tie_lo_T23Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y47__R0_BUF_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R0_INV_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y47__R1_BUF_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R1_INV_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R2_INV_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y47__R2_INV_1 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y47__R3_BUF_0 (.A(tie_lo_T23Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y48__R0_BUF_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R0_INV_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y48__R1_BUF_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R1_INV_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R2_INV_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y48__R2_INV_1 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y48__R3_BUF_0 (.A(tie_lo_T23Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y49__R0_BUF_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R0_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y49__R1_BUF_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R1_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R2_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y49__R2_INV_1 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y49__R3_BUF_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y4__R0_BUF_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R0_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y4__R1_BUF_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R1_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R2_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y4__R2_INV_1 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y4__R3_BUF_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y50__R0_BUF_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R0_INV_0 (.A(tie_lo_T23Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y50__R1_BUF_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R1_INV_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R2_INV_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y50__R2_INV_1 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y50__R3_BUF_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y51__R0_BUF_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R0_INV_0 (.A(tie_lo_T23Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y51__R1_BUF_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R1_INV_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R2_INV_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y51__R2_INV_1 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y51__R3_BUF_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y52__R0_BUF_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R0_INV_0 (.A(tie_lo_T23Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y52__R1_BUF_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R1_INV_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R2_INV_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y52__R2_INV_1 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y52__R3_BUF_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y53__R0_BUF_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R0_INV_0 (.A(tie_lo_T23Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y53__R1_BUF_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R1_INV_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R2_INV_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y53__R2_INV_1 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y53__R3_BUF_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y54__R0_BUF_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R0_INV_0 (.A(tie_lo_T23Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y54__R1_BUF_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R1_INV_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R2_INV_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y54__R2_INV_1 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y54__R3_BUF_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y55__R0_BUF_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R0_INV_0 (.A(tie_lo_T23Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y55__R1_BUF_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R1_INV_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R2_INV_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y55__R2_INV_1 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y55__R3_BUF_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y56__R0_BUF_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R0_INV_0 (.A(tie_lo_T23Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y56__R1_BUF_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R1_INV_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R2_INV_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y56__R2_INV_1 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y56__R3_BUF_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y57__R0_BUF_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R0_INV_0 (.A(tie_lo_T23Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y57__R1_BUF_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R1_INV_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R2_INV_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y57__R2_INV_1 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y57__R3_BUF_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y58__R0_BUF_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R0_INV_0 (.A(tie_lo_T23Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y58__R1_BUF_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R1_INV_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R2_INV_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y58__R2_INV_1 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y58__R3_BUF_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y59__R0_BUF_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R0_INV_0 (.A(tie_lo_T23Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y59__R1_BUF_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R1_INV_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R2_INV_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y59__R2_INV_1 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y59__R3_BUF_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y5__R0_BUF_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R0_INV_0 (.A(tie_lo_T23Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y5__R1_BUF_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R1_INV_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R2_INV_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y5__R2_INV_1 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y5__R3_BUF_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y60__R0_BUF_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R0_INV_0 (.A(tie_lo_T23Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y60__R1_BUF_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R1_INV_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R2_INV_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y60__R2_INV_1 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y60__R3_BUF_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y61__R0_BUF_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R0_INV_0 (.A(tie_lo_T23Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y61__R1_BUF_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R1_INV_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R2_INV_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y61__R2_INV_1 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y61__R3_BUF_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y62__R0_BUF_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R0_INV_0 (.A(tie_lo_T23Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y62__R1_BUF_0 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R1_INV_0 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R2_INV_0 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y62__R2_INV_1 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y62__R3_BUF_0 (.A(tie_lo_T23Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y63__R0_BUF_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R0_INV_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y63__R1_BUF_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R1_INV_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R2_INV_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y63__R2_INV_1 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y63__R3_BUF_0 (.A(tie_lo_T23Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y64__R0_BUF_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R0_INV_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y64__R1_BUF_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R1_INV_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R2_INV_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y64__R2_INV_1 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y64__R3_BUF_0 (.A(tie_lo_T23Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y65__R0_BUF_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R0_INV_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y65__R1_BUF_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R1_INV_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R2_INV_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y65__R2_INV_1 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y65__R3_BUF_0 (.A(tie_lo_T23Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y66__R0_BUF_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R0_INV_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y66__R1_BUF_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R1_INV_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R2_INV_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y66__R2_INV_1 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y66__R3_BUF_0 (.A(tie_lo_T23Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y67__R0_BUF_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R0_INV_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y67__R1_BUF_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R1_INV_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R2_INV_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y67__R2_INV_1 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y67__R3_BUF_0 (.A(tie_lo_T23Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y68__R0_BUF_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R0_INV_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y68__R1_BUF_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R1_INV_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R2_INV_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y68__R2_INV_1 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y68__R3_BUF_0 (.A(tie_lo_T23Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y69__R0_BUF_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R0_INV_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y69__R1_BUF_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R1_INV_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R2_INV_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y69__R2_INV_1 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y69__R3_BUF_0 (.A(tie_lo_T23Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y6__R0_BUF_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R0_INV_0 (.A(tie_lo_T23Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y6__R1_BUF_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R1_INV_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R2_INV_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y6__R2_INV_1 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y6__R3_BUF_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y70__R0_BUF_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R0_INV_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y70__R1_BUF_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R1_INV_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R2_INV_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y70__R2_INV_1 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y70__R3_BUF_0 (.A(tie_lo_T23Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y71__R0_BUF_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R0_INV_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y71__R1_BUF_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R1_INV_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R2_INV_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y71__R2_INV_1 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y71__R3_BUF_0 (.A(tie_lo_T23Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y72__R0_BUF_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R0_INV_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y72__R1_BUF_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R1_INV_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R2_INV_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y72__R2_INV_1 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y72__R3_BUF_0 (.A(tie_lo_T23Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y73__R0_BUF_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R0_INV_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y73__R1_BUF_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R1_INV_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R2_INV_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y73__R2_INV_1 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y73__R3_BUF_0 (.A(tie_lo_T23Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y74__R0_BUF_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R0_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y74__R1_BUF_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R1_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R2_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y74__R2_INV_1 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y74__R3_BUF_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y75__R0_BUF_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R0_INV_0 (.A(tie_lo_T23Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y75__R1_BUF_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R1_INV_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R2_INV_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y75__R2_INV_1 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y75__R3_BUF_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y76__R0_BUF_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R0_INV_0 (.A(tie_lo_T23Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y76__R1_BUF_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R1_INV_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R2_INV_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y76__R2_INV_1 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y76__R3_BUF_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y77__R0_BUF_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R0_INV_0 (.A(tie_lo_T23Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y77__R1_BUF_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R1_INV_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R2_INV_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y77__R2_INV_1 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y77__R3_BUF_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y78__R0_BUF_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R0_INV_0 (.A(tie_lo_T23Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y78__R1_BUF_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R1_INV_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R2_INV_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y78__R2_INV_1 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y78__R3_BUF_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y79__R0_BUF_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R0_INV_0 (.A(tie_lo_T23Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y79__R1_BUF_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R1_INV_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R2_INV_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y79__R2_INV_1 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y79__R3_BUF_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y7__R0_BUF_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R0_INV_0 (.A(tie_lo_T23Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y7__R1_BUF_0 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R1_INV_0 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R2_INV_0 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y7__R2_INV_1 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y7__R3_BUF_0 (.A(tie_lo_T23Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y80__R0_BUF_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R0_INV_0 (.A(tie_lo_T23Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y80__R1_BUF_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R1_INV_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R2_INV_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y80__R2_INV_1 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y80__R3_BUF_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y81__R0_BUF_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R0_INV_0 (.A(tie_lo_T23Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y81__R1_BUF_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R1_INV_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R2_INV_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y81__R2_INV_1 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y81__R3_BUF_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y82__R0_BUF_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R0_INV_0 (.A(tie_lo_T23Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y82__R1_BUF_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R1_INV_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R2_INV_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y82__R2_INV_1 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y82__R3_BUF_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y83__R0_BUF_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R0_INV_0 (.A(tie_lo_T23Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y83__R1_BUF_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R1_INV_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R2_INV_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y83__R2_INV_1 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y83__R3_BUF_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y84__R0_BUF_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R0_INV_0 (.A(tie_lo_T23Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y84__R1_BUF_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R1_INV_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R2_INV_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y84__R2_INV_1 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y84__R3_BUF_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y85__R0_BUF_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R0_INV_0 (.A(tie_lo_T23Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y85__R1_BUF_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R1_INV_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R2_INV_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y85__R2_INV_1 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y85__R3_BUF_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y86__R0_BUF_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R0_INV_0 (.A(tie_lo_T23Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y86__R1_BUF_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R1_INV_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R2_INV_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y86__R2_INV_1 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y86__R3_BUF_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y87__R0_BUF_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R0_INV_0 (.A(tie_lo_T23Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y87__R1_BUF_0 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R1_INV_0 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R2_INV_0 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y87__R2_INV_1 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y87__R3_BUF_0 (.A(tie_lo_T23Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y88__R0_BUF_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R0_INV_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y88__R1_BUF_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R1_INV_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R2_INV_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y88__R2_INV_1 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y88__R3_BUF_0 (.A(tie_lo_T23Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y89__R0_BUF_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R0_INV_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y89__R1_BUF_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R1_INV_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R2_INV_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y89__R2_INV_1 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y89__R3_BUF_0 (.A(tie_lo_T23Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y8__R0_BUF_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R0_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y8__R1_BUF_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R1_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R2_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y8__R2_INV_1 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y8__R3_BUF_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y9__R0_BUF_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R0_INV_0 (.A(tie_lo_T23Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y9__R1_BUF_0 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R1_INV_0 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T23Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R2_INV_0 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T23Y9__R2_INV_1 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T23Y9__R3_BUF_0 (.A(tie_lo_T23Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y0__R0_BUF_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R0_INV_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y0__R1_BUF_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R1_INV_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R2_INV_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y0__R2_INV_1 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y0__R3_BUF_0 (.A(tie_lo_T24Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y10__R0_BUF_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R0_INV_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y10__R1_BUF_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R1_INV_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R2_INV_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y10__R2_INV_1 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y10__R3_BUF_0 (.A(tie_lo_T24Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y11__R0_BUF_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R0_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y11__R1_BUF_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R1_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R2_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y11__R2_INV_1 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y11__R3_BUF_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y12__R0_BUF_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R0_INV_0 (.A(tie_lo_T24Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y12__R1_BUF_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R1_INV_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R2_INV_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y12__R2_INV_1 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y12__R3_BUF_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y13__R0_BUF_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R0_INV_0 (.A(tie_lo_T24Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y13__R1_BUF_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R1_INV_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R2_INV_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y13__R2_INV_1 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y13__R3_BUF_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y14__R0_BUF_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R0_INV_0 (.A(tie_lo_T24Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y14__R1_BUF_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R1_INV_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R2_INV_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y14__R2_INV_1 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y14__R3_BUF_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y15__R0_BUF_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R0_INV_0 (.A(tie_lo_T24Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y15__R1_BUF_0 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R1_INV_0 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R2_INV_0 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y15__R2_INV_1 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y15__R3_BUF_0 (.A(tie_lo_T24Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y16__R0_BUF_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R0_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y16__R1_BUF_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R1_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R2_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y16__R2_INV_1 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y16__R3_BUF_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y17__R0_BUF_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R0_INV_0 (.A(tie_lo_T24Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y17__R1_BUF_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R1_INV_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R2_INV_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y17__R2_INV_1 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y17__R3_BUF_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y18__R0_BUF_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R0_INV_0 (.A(tie_lo_T24Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y18__R1_BUF_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R1_INV_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R2_INV_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y18__R2_INV_1 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y18__R3_BUF_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y19__R0_BUF_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R0_INV_0 (.A(tie_lo_T24Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y19__R1_BUF_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R1_INV_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R2_INV_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y19__R2_INV_1 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y19__R3_BUF_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y1__R0_BUF_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R0_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y1__R1_BUF_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R1_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R2_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y1__R2_INV_1 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y1__R3_BUF_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y20__R0_BUF_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R0_INV_0 (.A(tie_lo_T24Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y20__R1_BUF_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R1_INV_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R2_INV_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y20__R2_INV_1 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y20__R3_BUF_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y21__R0_BUF_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R0_INV_0 (.A(tie_lo_T24Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y21__R1_BUF_0 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R1_INV_0 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R2_INV_0 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y21__R2_INV_1 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y21__R3_BUF_0 (.A(tie_lo_T24Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y22__R0_BUF_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R0_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y22__R1_BUF_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R1_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R2_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y22__R2_INV_1 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y22__R3_BUF_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y23__R0_BUF_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R0_INV_0 (.A(tie_lo_T24Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y23__R1_BUF_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R1_INV_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R2_INV_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y23__R2_INV_1 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y23__R3_BUF_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y24__R0_BUF_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R0_INV_0 (.A(tie_lo_T24Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y24__R1_BUF_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R1_INV_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R2_INV_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y24__R2_INV_1 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y24__R3_BUF_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y25__R0_BUF_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R0_INV_0 (.A(tie_lo_T24Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y25__R1_BUF_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R1_INV_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R2_INV_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y25__R2_INV_1 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y25__R3_BUF_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y26__R0_BUF_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R0_INV_0 (.A(tie_lo_T24Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y26__R1_BUF_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R1_INV_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R2_INV_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y26__R2_INV_1 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y26__R3_BUF_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y27__R0_BUF_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R0_INV_0 (.A(tie_lo_T24Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y27__R1_BUF_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R1_INV_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R2_INV_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y27__R2_INV_1 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y27__R3_BUF_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y28__R0_BUF_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R0_INV_0 (.A(tie_lo_T24Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y28__R1_BUF_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R1_INV_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R2_INV_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y28__R2_INV_1 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y28__R3_BUF_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y29__R0_BUF_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R0_INV_0 (.A(tie_lo_T24Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y29__R1_BUF_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R1_INV_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R2_INV_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y29__R2_INV_1 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y29__R3_BUF_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y2__R0_BUF_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R0_INV_0 (.A(tie_lo_T24Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y2__R1_BUF_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R1_INV_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R2_INV_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y2__R2_INV_1 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y2__R3_BUF_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y30__R0_BUF_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R0_INV_0 (.A(tie_lo_T24Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y30__R1_BUF_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R1_INV_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R2_INV_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y30__R2_INV_1 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y30__R3_BUF_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y31__R0_BUF_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R0_INV_0 (.A(tie_lo_T24Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y31__R1_BUF_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R1_INV_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R2_INV_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y31__R2_INV_1 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y31__R3_BUF_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y32__R0_BUF_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R0_INV_0 (.A(tie_lo_T24Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y32__R1_BUF_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R1_INV_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R2_INV_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y32__R2_INV_1 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y32__R3_BUF_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y33__R0_BUF_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R0_INV_0 (.A(tie_lo_T24Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y33__R1_BUF_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R1_INV_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R2_INV_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y33__R2_INV_1 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y33__R3_BUF_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y34__R0_BUF_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R0_INV_0 (.A(tie_lo_T24Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y34__R1_BUF_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R1_INV_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R2_INV_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y34__R2_INV_1 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y34__R3_BUF_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y35__R0_BUF_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R0_INV_0 (.A(tie_lo_T24Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y35__R1_BUF_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R1_INV_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R2_INV_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y35__R2_INV_1 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y35__R3_BUF_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y36__R0_BUF_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R0_INV_0 (.A(tie_lo_T24Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y36__R1_BUF_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R1_INV_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R2_INV_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y36__R2_INV_1 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y36__R3_BUF_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y37__R0_BUF_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R0_INV_0 (.A(tie_lo_T24Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y37__R1_BUF_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R1_INV_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R2_INV_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y37__R2_INV_1 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y37__R3_BUF_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y38__R0_BUF_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R0_INV_0 (.A(tie_lo_T24Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y38__R1_BUF_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R1_INV_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R2_INV_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y38__R2_INV_1 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y38__R3_BUF_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y39__R0_BUF_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R0_INV_0 (.A(tie_lo_T24Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y39__R1_BUF_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R1_INV_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R2_INV_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y39__R2_INV_1 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y39__R3_BUF_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y3__R0_BUF_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R0_INV_0 (.A(tie_lo_T24Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y3__R1_BUF_0 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R1_INV_0 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R2_INV_0 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y3__R2_INV_1 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y3__R3_BUF_0 (.A(tie_lo_T24Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y40__R0_BUF_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R0_INV_0 (.A(tie_lo_T24Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y40__R1_BUF_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R1_INV_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R2_INV_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y40__R2_INV_1 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y40__R3_BUF_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y41__R0_BUF_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R0_INV_0 (.A(tie_lo_T24Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y41__R1_BUF_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R1_INV_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R2_INV_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y41__R2_INV_1 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y41__R3_BUF_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y42__R0_BUF_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R0_INV_0 (.A(tie_lo_T24Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y42__R1_BUF_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R1_INV_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R2_INV_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y42__R2_INV_1 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y42__R3_BUF_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y43__R0_BUF_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R0_INV_0 (.A(tie_lo_T24Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y43__R1_BUF_0 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R1_INV_0 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R2_INV_0 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y43__R2_INV_1 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y43__R3_BUF_0 (.A(tie_lo_T24Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y44__R0_BUF_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R0_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y44__R1_BUF_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R1_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R2_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y44__R2_INV_1 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y44__R3_BUF_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y45__R0_BUF_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R0_INV_0 (.A(tie_lo_T24Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y45__R1_BUF_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R1_INV_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R2_INV_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y45__R2_INV_1 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y45__R3_BUF_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y46__R0_BUF_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R0_INV_0 (.A(tie_lo_T24Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y46__R1_BUF_0 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R1_INV_0 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R2_INV_0 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y46__R2_INV_1 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y46__R3_BUF_0 (.A(tie_lo_T24Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y47__R0_BUF_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R0_INV_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y47__R1_BUF_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R1_INV_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R2_INV_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y47__R2_INV_1 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y47__R3_BUF_0 (.A(tie_lo_T24Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y48__R0_BUF_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R0_INV_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y48__R1_BUF_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R1_INV_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R2_INV_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y48__R2_INV_1 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y48__R3_BUF_0 (.A(tie_lo_T24Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y49__R0_BUF_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R0_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y49__R1_BUF_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R1_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R2_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y49__R2_INV_1 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y49__R3_BUF_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y4__R0_BUF_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R0_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y4__R1_BUF_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R1_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R2_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y4__R2_INV_1 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y4__R3_BUF_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y50__R0_BUF_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R0_INV_0 (.A(tie_lo_T24Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y50__R1_BUF_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R1_INV_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R2_INV_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y50__R2_INV_1 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y50__R3_BUF_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y51__R0_BUF_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R0_INV_0 (.A(tie_lo_T24Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y51__R1_BUF_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R1_INV_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R2_INV_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y51__R2_INV_1 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y51__R3_BUF_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y52__R0_BUF_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R0_INV_0 (.A(tie_lo_T24Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y52__R1_BUF_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R1_INV_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R2_INV_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y52__R2_INV_1 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y52__R3_BUF_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y53__R0_BUF_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R0_INV_0 (.A(tie_lo_T24Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y53__R1_BUF_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R1_INV_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R2_INV_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y53__R2_INV_1 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y53__R3_BUF_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y54__R0_BUF_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R0_INV_0 (.A(tie_lo_T24Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y54__R1_BUF_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R1_INV_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R2_INV_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y54__R2_INV_1 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y54__R3_BUF_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y55__R0_BUF_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R0_INV_0 (.A(tie_lo_T24Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y55__R1_BUF_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R1_INV_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R2_INV_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y55__R2_INV_1 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y55__R3_BUF_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y56__R0_BUF_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R0_INV_0 (.A(tie_lo_T24Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y56__R1_BUF_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R1_INV_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R2_INV_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y56__R2_INV_1 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y56__R3_BUF_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y57__R0_BUF_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R0_INV_0 (.A(tie_lo_T24Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y57__R1_BUF_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R1_INV_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R2_INV_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y57__R2_INV_1 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y57__R3_BUF_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y58__R0_BUF_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R0_INV_0 (.A(tie_lo_T24Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y58__R1_BUF_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R1_INV_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R2_INV_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y58__R2_INV_1 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y58__R3_BUF_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y59__R0_BUF_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R0_INV_0 (.A(tie_lo_T24Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y59__R1_BUF_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R1_INV_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R2_INV_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y59__R2_INV_1 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y59__R3_BUF_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y5__R0_BUF_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R0_INV_0 (.A(tie_lo_T24Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y5__R1_BUF_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R1_INV_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R2_INV_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y5__R2_INV_1 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y5__R3_BUF_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y60__R0_BUF_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R0_INV_0 (.A(tie_lo_T24Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y60__R1_BUF_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R1_INV_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R2_INV_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y60__R2_INV_1 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y60__R3_BUF_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y61__R0_BUF_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R0_INV_0 (.A(tie_lo_T24Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y61__R1_BUF_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R1_INV_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R2_INV_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y61__R2_INV_1 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y61__R3_BUF_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y62__R0_BUF_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R0_INV_0 (.A(tie_lo_T24Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y62__R1_BUF_0 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R1_INV_0 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R2_INV_0 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y62__R2_INV_1 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y62__R3_BUF_0 (.A(tie_lo_T24Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y63__R0_BUF_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R0_INV_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y63__R1_BUF_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R1_INV_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R2_INV_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y63__R2_INV_1 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y63__R3_BUF_0 (.A(tie_lo_T24Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y64__R0_BUF_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R0_INV_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y64__R1_BUF_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R1_INV_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R2_INV_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y64__R2_INV_1 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y64__R3_BUF_0 (.A(tie_lo_T24Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y65__R0_BUF_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R0_INV_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y65__R1_BUF_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R1_INV_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R2_INV_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y65__R2_INV_1 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y65__R3_BUF_0 (.A(tie_lo_T24Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y66__R0_BUF_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R0_INV_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y66__R1_BUF_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R1_INV_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R2_INV_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y66__R2_INV_1 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y66__R3_BUF_0 (.A(tie_lo_T24Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y67__R0_BUF_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R0_INV_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y67__R1_BUF_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R1_INV_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R2_INV_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y67__R2_INV_1 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y67__R3_BUF_0 (.A(tie_lo_T24Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y68__R0_BUF_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R0_INV_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y68__R1_BUF_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R1_INV_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R2_INV_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y68__R2_INV_1 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y68__R3_BUF_0 (.A(tie_lo_T24Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y69__R0_BUF_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R0_INV_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y69__R1_BUF_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R1_INV_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R2_INV_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y69__R2_INV_1 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y69__R3_BUF_0 (.A(tie_lo_T24Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y6__R0_BUF_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R0_INV_0 (.A(tie_lo_T24Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y6__R1_BUF_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R1_INV_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R2_INV_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y6__R2_INV_1 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y6__R3_BUF_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y70__R0_BUF_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R0_INV_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y70__R1_BUF_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R1_INV_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R2_INV_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y70__R2_INV_1 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y70__R3_BUF_0 (.A(tie_lo_T24Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y71__R0_BUF_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R0_INV_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y71__R1_BUF_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R1_INV_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R2_INV_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y71__R2_INV_1 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y71__R3_BUF_0 (.A(tie_lo_T24Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y72__R0_BUF_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R0_INV_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y72__R1_BUF_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R1_INV_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R2_INV_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y72__R2_INV_1 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y72__R3_BUF_0 (.A(tie_lo_T24Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y73__R0_BUF_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R0_INV_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y73__R1_BUF_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R1_INV_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R2_INV_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y73__R2_INV_1 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y73__R3_BUF_0 (.A(tie_lo_T24Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y74__R0_BUF_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R0_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y74__R1_BUF_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R1_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R2_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y74__R2_INV_1 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y74__R3_BUF_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y75__R0_BUF_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R0_INV_0 (.A(tie_lo_T24Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y75__R1_BUF_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R1_INV_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R2_INV_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y75__R2_INV_1 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y75__R3_BUF_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y76__R0_BUF_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R0_INV_0 (.A(tie_lo_T24Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y76__R1_BUF_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R1_INV_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R2_INV_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y76__R2_INV_1 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y76__R3_BUF_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y77__R0_BUF_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R0_INV_0 (.A(tie_lo_T24Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y77__R1_BUF_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R1_INV_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R2_INV_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y77__R2_INV_1 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y77__R3_BUF_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y78__R0_BUF_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R0_INV_0 (.A(tie_lo_T24Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y78__R1_BUF_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R1_INV_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R2_INV_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y78__R2_INV_1 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y78__R3_BUF_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y79__R0_BUF_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R0_INV_0 (.A(tie_lo_T24Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y79__R1_BUF_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R1_INV_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R2_INV_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y79__R2_INV_1 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y79__R3_BUF_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y7__R0_BUF_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R0_INV_0 (.A(tie_lo_T24Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y7__R1_BUF_0 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R1_INV_0 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R2_INV_0 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y7__R2_INV_1 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y7__R3_BUF_0 (.A(tie_lo_T24Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y80__R0_BUF_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R0_INV_0 (.A(tie_lo_T24Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y80__R1_BUF_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R1_INV_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R2_INV_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y80__R2_INV_1 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y80__R3_BUF_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y81__R0_BUF_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R0_INV_0 (.A(tie_lo_T24Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y81__R1_BUF_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R1_INV_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R2_INV_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y81__R2_INV_1 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y81__R3_BUF_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y82__R0_BUF_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R0_INV_0 (.A(tie_lo_T24Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y82__R1_BUF_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R1_INV_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R2_INV_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y82__R2_INV_1 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y82__R3_BUF_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y83__R0_BUF_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R0_INV_0 (.A(tie_lo_T24Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y83__R1_BUF_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R1_INV_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R2_INV_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y83__R2_INV_1 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y83__R3_BUF_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y84__R0_BUF_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R0_INV_0 (.A(tie_lo_T24Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y84__R1_BUF_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R1_INV_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R2_INV_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y84__R2_INV_1 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y84__R3_BUF_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y85__R0_BUF_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R0_INV_0 (.A(tie_lo_T24Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y85__R1_BUF_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R1_INV_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R2_INV_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y85__R2_INV_1 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y85__R3_BUF_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y86__R0_BUF_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R0_INV_0 (.A(tie_lo_T24Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y86__R1_BUF_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R1_INV_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R2_INV_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y86__R2_INV_1 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y86__R3_BUF_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y87__R0_BUF_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R0_INV_0 (.A(tie_lo_T24Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y87__R1_BUF_0 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R1_INV_0 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R2_INV_0 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y87__R2_INV_1 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y87__R3_BUF_0 (.A(tie_lo_T24Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y88__R0_BUF_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R0_INV_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y88__R1_BUF_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R1_INV_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R2_INV_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y88__R2_INV_1 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y88__R3_BUF_0 (.A(tie_lo_T24Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y89__R0_BUF_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R0_INV_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y89__R1_BUF_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R1_INV_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R2_INV_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y89__R2_INV_1 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y89__R3_BUF_0 (.A(tie_lo_T24Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y8__R0_BUF_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R0_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y8__R1_BUF_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R1_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R2_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y8__R2_INV_1 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y8__R3_BUF_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y9__R0_BUF_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R0_INV_0 (.A(tie_lo_T24Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y9__R1_BUF_0 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R1_INV_0 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T24Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R2_INV_0 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T24Y9__R2_INV_1 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T24Y9__R3_BUF_0 (.A(tie_lo_T24Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y0__R0_BUF_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R0_INV_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y0__R1_BUF_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R1_INV_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R2_INV_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y0__R2_INV_1 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y0__R3_BUF_0 (.A(tie_lo_T25Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y10__R0_BUF_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R0_INV_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y10__R1_BUF_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R1_INV_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R2_INV_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y10__R2_INV_1 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y10__R3_BUF_0 (.A(tie_lo_T25Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y11__R0_BUF_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R0_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y11__R1_BUF_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R1_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R2_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y11__R2_INV_1 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y11__R3_BUF_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y12__R0_BUF_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R0_INV_0 (.A(tie_lo_T25Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y12__R1_BUF_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R1_INV_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R2_INV_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y12__R2_INV_1 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y12__R3_BUF_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y13__R0_BUF_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R0_INV_0 (.A(tie_lo_T25Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y13__R1_BUF_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R1_INV_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R2_INV_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y13__R2_INV_1 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y13__R3_BUF_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y14__R0_BUF_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R0_INV_0 (.A(tie_lo_T25Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y14__R1_BUF_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R1_INV_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R2_INV_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y14__R2_INV_1 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y14__R3_BUF_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y15__R0_BUF_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R0_INV_0 (.A(tie_lo_T25Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y15__R1_BUF_0 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R1_INV_0 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R2_INV_0 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y15__R2_INV_1 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y15__R3_BUF_0 (.A(tie_lo_T25Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y16__R0_BUF_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R0_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y16__R1_BUF_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R1_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R2_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y16__R2_INV_1 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y16__R3_BUF_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y17__R0_BUF_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R0_INV_0 (.A(tie_lo_T25Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y17__R1_BUF_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R1_INV_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R2_INV_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y17__R2_INV_1 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y17__R3_BUF_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y18__R0_BUF_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R0_INV_0 (.A(tie_lo_T25Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y18__R1_BUF_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R1_INV_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R2_INV_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y18__R2_INV_1 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y18__R3_BUF_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y19__R0_BUF_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R0_INV_0 (.A(tie_lo_T25Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y19__R1_BUF_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R1_INV_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R2_INV_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y19__R2_INV_1 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y19__R3_BUF_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y1__R0_BUF_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R0_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y1__R1_BUF_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R1_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R2_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y1__R2_INV_1 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y1__R3_BUF_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y20__R0_BUF_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R0_INV_0 (.A(tie_lo_T25Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y20__R1_BUF_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R1_INV_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R2_INV_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y20__R2_INV_1 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y20__R3_BUF_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y21__R0_BUF_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R0_INV_0 (.A(tie_lo_T25Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y21__R1_BUF_0 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R1_INV_0 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R2_INV_0 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y21__R2_INV_1 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y21__R3_BUF_0 (.A(tie_lo_T25Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y22__R0_BUF_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R0_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y22__R1_BUF_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R1_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R2_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y22__R2_INV_1 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y22__R3_BUF_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y23__R0_BUF_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R0_INV_0 (.A(tie_lo_T25Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y23__R1_BUF_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R1_INV_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R2_INV_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y23__R2_INV_1 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y23__R3_BUF_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y24__R0_BUF_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R0_INV_0 (.A(tie_lo_T25Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y24__R1_BUF_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R1_INV_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R2_INV_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y24__R2_INV_1 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y24__R3_BUF_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y25__R0_BUF_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R0_INV_0 (.A(tie_lo_T25Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y25__R1_BUF_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R1_INV_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R2_INV_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y25__R2_INV_1 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y25__R3_BUF_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y26__R0_BUF_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R0_INV_0 (.A(tie_lo_T25Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y26__R1_BUF_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R1_INV_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R2_INV_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y26__R2_INV_1 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y26__R3_BUF_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y27__R0_BUF_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R0_INV_0 (.A(tie_lo_T25Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y27__R1_BUF_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R1_INV_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R2_INV_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y27__R2_INV_1 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y27__R3_BUF_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y28__R0_BUF_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R0_INV_0 (.A(tie_lo_T25Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y28__R1_BUF_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R1_INV_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R2_INV_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y28__R2_INV_1 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y28__R3_BUF_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y29__R0_BUF_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R0_INV_0 (.A(tie_lo_T25Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y29__R1_BUF_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R1_INV_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R2_INV_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y29__R2_INV_1 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y29__R3_BUF_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y2__R0_BUF_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R0_INV_0 (.A(tie_lo_T25Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y2__R1_BUF_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R1_INV_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R2_INV_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y2__R2_INV_1 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y2__R3_BUF_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y30__R0_BUF_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R0_INV_0 (.A(tie_lo_T25Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y30__R1_BUF_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R1_INV_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R2_INV_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y30__R2_INV_1 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y30__R3_BUF_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y31__R0_BUF_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R0_INV_0 (.A(tie_lo_T25Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y31__R1_BUF_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R1_INV_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R2_INV_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y31__R2_INV_1 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y31__R3_BUF_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y32__R0_BUF_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R0_INV_0 (.A(tie_lo_T25Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y32__R1_BUF_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R1_INV_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R2_INV_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y32__R2_INV_1 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y32__R3_BUF_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y33__R0_BUF_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R0_INV_0 (.A(tie_lo_T25Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y33__R1_BUF_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R1_INV_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R2_INV_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y33__R2_INV_1 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y33__R3_BUF_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y34__R0_BUF_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R0_INV_0 (.A(tie_lo_T25Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y34__R1_BUF_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R1_INV_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R2_INV_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y34__R2_INV_1 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y34__R3_BUF_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y35__R0_BUF_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R0_INV_0 (.A(tie_lo_T25Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y35__R1_BUF_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R1_INV_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R2_INV_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y35__R2_INV_1 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y35__R3_BUF_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y36__R0_BUF_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R0_INV_0 (.A(tie_lo_T25Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y36__R1_BUF_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R1_INV_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R2_INV_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y36__R2_INV_1 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y36__R3_BUF_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y37__R0_BUF_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R0_INV_0 (.A(tie_lo_T25Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y37__R1_BUF_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R1_INV_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R2_INV_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y37__R2_INV_1 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y37__R3_BUF_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y38__R0_BUF_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R0_INV_0 (.A(tie_lo_T25Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y38__R1_BUF_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R1_INV_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R2_INV_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y38__R2_INV_1 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y38__R3_BUF_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y39__R0_BUF_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R0_INV_0 (.A(tie_lo_T25Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y39__R1_BUF_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R1_INV_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R2_INV_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y39__R2_INV_1 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y39__R3_BUF_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y3__R0_BUF_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R0_INV_0 (.A(tie_lo_T25Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y3__R1_BUF_0 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R1_INV_0 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R2_INV_0 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y3__R2_INV_1 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y3__R3_BUF_0 (.A(tie_lo_T25Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y40__R0_BUF_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R0_INV_0 (.A(tie_lo_T25Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y40__R1_BUF_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R1_INV_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R2_INV_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y40__R2_INV_1 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y40__R3_BUF_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y41__R0_BUF_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R0_INV_0 (.A(tie_lo_T25Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y41__R1_BUF_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R1_INV_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R2_INV_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y41__R2_INV_1 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y41__R3_BUF_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y42__R0_BUF_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R0_INV_0 (.A(tie_lo_T25Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y42__R1_BUF_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R1_INV_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R2_INV_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y42__R2_INV_1 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y42__R3_BUF_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y43__R0_BUF_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R0_INV_0 (.A(tie_lo_T25Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y43__R1_BUF_0 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R1_INV_0 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R2_INV_0 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y43__R2_INV_1 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y43__R3_BUF_0 (.A(tie_lo_T25Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y44__R0_BUF_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R0_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y44__R1_BUF_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R1_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R2_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y44__R2_INV_1 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y44__R3_BUF_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y45__R0_BUF_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R0_INV_0 (.A(tie_lo_T25Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y45__R1_BUF_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R1_INV_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R2_INV_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y45__R2_INV_1 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y45__R3_BUF_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y46__R0_BUF_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R0_INV_0 (.A(tie_lo_T25Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y46__R1_BUF_0 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R1_INV_0 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R2_INV_0 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y46__R2_INV_1 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y46__R3_BUF_0 (.A(tie_lo_T25Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y47__R0_BUF_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R0_INV_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y47__R1_BUF_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R1_INV_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R2_INV_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y47__R2_INV_1 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y47__R3_BUF_0 (.A(tie_lo_T25Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y48__R0_BUF_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R0_INV_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y48__R1_BUF_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R1_INV_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R2_INV_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y48__R2_INV_1 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y48__R3_BUF_0 (.A(tie_lo_T25Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y49__R0_BUF_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R0_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y49__R1_BUF_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R1_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R2_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y49__R2_INV_1 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y49__R3_BUF_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y4__R0_BUF_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R0_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y4__R1_BUF_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R1_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R2_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y4__R2_INV_1 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y4__R3_BUF_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y50__R0_BUF_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R0_INV_0 (.A(tie_lo_T25Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y50__R1_BUF_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R1_INV_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R2_INV_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y50__R2_INV_1 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y50__R3_BUF_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y51__R0_BUF_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R0_INV_0 (.A(tie_lo_T25Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y51__R1_BUF_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R1_INV_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R2_INV_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y51__R2_INV_1 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y51__R3_BUF_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y52__R0_BUF_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R0_INV_0 (.A(tie_lo_T25Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y52__R1_BUF_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R1_INV_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R2_INV_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y52__R2_INV_1 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y52__R3_BUF_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y53__R0_BUF_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R0_INV_0 (.A(tie_lo_T25Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y53__R1_BUF_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R1_INV_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R2_INV_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y53__R2_INV_1 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y53__R3_BUF_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y54__R0_BUF_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R0_INV_0 (.A(tie_lo_T25Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y54__R1_BUF_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R1_INV_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R2_INV_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y54__R2_INV_1 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y54__R3_BUF_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y55__R0_BUF_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R0_INV_0 (.A(tie_lo_T25Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y55__R1_BUF_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R1_INV_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R2_INV_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y55__R2_INV_1 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y55__R3_BUF_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y56__R0_BUF_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R0_INV_0 (.A(tie_lo_T25Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y56__R1_BUF_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R1_INV_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R2_INV_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y56__R2_INV_1 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y56__R3_BUF_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y57__R0_BUF_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R0_INV_0 (.A(tie_lo_T25Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y57__R1_BUF_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R1_INV_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R2_INV_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y57__R2_INV_1 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y57__R3_BUF_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y58__R0_BUF_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R0_INV_0 (.A(tie_lo_T25Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y58__R1_BUF_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R1_INV_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R2_INV_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y58__R2_INV_1 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y58__R3_BUF_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y59__R0_BUF_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R0_INV_0 (.A(tie_lo_T25Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y59__R1_BUF_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R1_INV_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R2_INV_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y59__R2_INV_1 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y59__R3_BUF_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y5__R0_BUF_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R0_INV_0 (.A(tie_lo_T25Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y5__R1_BUF_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R1_INV_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R2_INV_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y5__R2_INV_1 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y5__R3_BUF_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y60__R0_BUF_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R0_INV_0 (.A(tie_lo_T25Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y60__R1_BUF_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R1_INV_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R2_INV_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y60__R2_INV_1 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y60__R3_BUF_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y61__R0_BUF_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R0_INV_0 (.A(tie_lo_T25Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y61__R1_BUF_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R1_INV_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R2_INV_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y61__R2_INV_1 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y61__R3_BUF_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y62__R0_BUF_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R0_INV_0 (.A(tie_lo_T25Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y62__R1_BUF_0 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R1_INV_0 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R2_INV_0 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y62__R2_INV_1 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y62__R3_BUF_0 (.A(tie_lo_T25Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y63__R0_BUF_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R0_INV_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y63__R1_BUF_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R1_INV_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R2_INV_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y63__R2_INV_1 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y63__R3_BUF_0 (.A(tie_lo_T25Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y64__R0_BUF_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R0_INV_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y64__R1_BUF_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R1_INV_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R2_INV_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y64__R2_INV_1 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y64__R3_BUF_0 (.A(tie_lo_T25Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y65__R0_BUF_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R0_INV_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y65__R1_BUF_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R1_INV_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R2_INV_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y65__R2_INV_1 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y65__R3_BUF_0 (.A(tie_lo_T25Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y66__R0_BUF_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R0_INV_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y66__R1_BUF_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R1_INV_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R2_INV_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y66__R2_INV_1 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y66__R3_BUF_0 (.A(tie_lo_T25Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y67__R0_BUF_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R0_INV_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y67__R1_BUF_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R1_INV_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R2_INV_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y67__R2_INV_1 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y67__R3_BUF_0 (.A(tie_lo_T25Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y68__R0_BUF_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R0_INV_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y68__R1_BUF_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R1_INV_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R2_INV_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y68__R2_INV_1 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y68__R3_BUF_0 (.A(tie_lo_T25Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y69__R0_BUF_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R0_INV_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y69__R1_BUF_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R1_INV_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R2_INV_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y69__R2_INV_1 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y69__R3_BUF_0 (.A(tie_lo_T25Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y6__R0_BUF_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R0_INV_0 (.A(tie_lo_T25Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y6__R1_BUF_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R1_INV_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R2_INV_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y6__R2_INV_1 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y6__R3_BUF_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y70__R0_BUF_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R0_INV_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y70__R1_BUF_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R1_INV_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R2_INV_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y70__R2_INV_1 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y70__R3_BUF_0 (.A(tie_lo_T25Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y71__R0_BUF_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R0_INV_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y71__R1_BUF_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R1_INV_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R2_INV_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y71__R2_INV_1 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y71__R3_BUF_0 (.A(tie_lo_T25Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y72__R0_BUF_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R0_INV_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y72__R1_BUF_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R1_INV_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R2_INV_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y72__R2_INV_1 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y72__R3_BUF_0 (.A(tie_lo_T25Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y73__R0_BUF_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R0_INV_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y73__R1_BUF_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R1_INV_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R2_INV_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y73__R2_INV_1 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y73__R3_BUF_0 (.A(tie_lo_T25Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y74__R0_BUF_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R0_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y74__R1_BUF_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R1_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R2_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y74__R2_INV_1 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y74__R3_BUF_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y75__R0_BUF_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R0_INV_0 (.A(tie_lo_T25Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y75__R1_BUF_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R1_INV_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R2_INV_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y75__R2_INV_1 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y75__R3_BUF_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y76__R0_BUF_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R0_INV_0 (.A(tie_lo_T25Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y76__R1_BUF_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R1_INV_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R2_INV_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y76__R2_INV_1 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y76__R3_BUF_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y77__R0_BUF_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R0_INV_0 (.A(tie_lo_T25Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y77__R1_BUF_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R1_INV_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R2_INV_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y77__R2_INV_1 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y77__R3_BUF_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y78__R0_BUF_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R0_INV_0 (.A(tie_lo_T25Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y78__R1_BUF_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R1_INV_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R2_INV_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y78__R2_INV_1 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y78__R3_BUF_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y79__R0_BUF_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R0_INV_0 (.A(tie_lo_T25Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y79__R1_BUF_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R1_INV_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R2_INV_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y79__R2_INV_1 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y79__R3_BUF_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y7__R0_BUF_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R0_INV_0 (.A(tie_lo_T25Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y7__R1_BUF_0 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R1_INV_0 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R2_INV_0 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y7__R2_INV_1 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y7__R3_BUF_0 (.A(tie_lo_T25Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y80__R0_BUF_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R0_INV_0 (.A(tie_lo_T25Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y80__R1_BUF_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R1_INV_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R2_INV_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y80__R2_INV_1 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y80__R3_BUF_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y81__R0_BUF_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R0_INV_0 (.A(tie_lo_T25Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y81__R1_BUF_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R1_INV_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R2_INV_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y81__R2_INV_1 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y81__R3_BUF_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y82__R0_BUF_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R0_INV_0 (.A(tie_lo_T25Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y82__R1_BUF_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R1_INV_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R2_INV_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y82__R2_INV_1 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y82__R3_BUF_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y83__R0_BUF_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R0_INV_0 (.A(tie_lo_T25Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y83__R1_BUF_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R1_INV_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R2_INV_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y83__R2_INV_1 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y83__R3_BUF_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y84__R0_BUF_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R0_INV_0 (.A(tie_lo_T25Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y84__R1_BUF_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R1_INV_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R2_INV_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y84__R2_INV_1 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y84__R3_BUF_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y85__R0_BUF_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R0_INV_0 (.A(tie_lo_T25Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y85__R1_BUF_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R1_INV_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R2_INV_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y85__R2_INV_1 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y85__R3_BUF_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y86__R0_BUF_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R0_INV_0 (.A(tie_lo_T25Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y86__R1_BUF_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R1_INV_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R2_INV_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y86__R2_INV_1 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y86__R3_BUF_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y87__R0_BUF_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R0_INV_0 (.A(tie_lo_T25Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y87__R1_BUF_0 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R1_INV_0 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R2_INV_0 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y87__R2_INV_1 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y87__R3_BUF_0 (.A(tie_lo_T25Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y88__R0_BUF_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R0_INV_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y88__R1_BUF_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R1_INV_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R2_INV_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y88__R2_INV_1 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y88__R3_BUF_0 (.A(tie_lo_T25Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y89__R0_BUF_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R0_INV_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y89__R1_BUF_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R1_INV_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R2_INV_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y89__R2_INV_1 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y89__R3_BUF_0 (.A(tie_lo_T25Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y8__R0_BUF_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R0_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y8__R1_BUF_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R1_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R2_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y8__R2_INV_1 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y8__R3_BUF_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y9__R0_BUF_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R0_INV_0 (.A(tie_lo_T25Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y9__R1_BUF_0 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R1_INV_0 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T25Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R2_INV_0 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T25Y9__R2_INV_1 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T25Y9__R3_BUF_0 (.A(tie_lo_T25Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y0__R0_BUF_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R0_INV_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y0__R1_BUF_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R1_INV_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R2_INV_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y0__R2_INV_1 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y0__R3_BUF_0 (.A(tie_lo_T26Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y10__R0_BUF_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R0_INV_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y10__R1_BUF_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R1_INV_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R2_INV_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y10__R2_INV_1 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y10__R3_BUF_0 (.A(tie_lo_T26Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y11__R0_BUF_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R0_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y11__R1_BUF_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R1_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R2_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y11__R2_INV_1 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y11__R3_BUF_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y12__R0_BUF_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R0_INV_0 (.A(tie_lo_T26Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y12__R1_BUF_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R1_INV_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R2_INV_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y12__R2_INV_1 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y12__R3_BUF_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y13__R0_BUF_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R0_INV_0 (.A(tie_lo_T26Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y13__R1_BUF_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R1_INV_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R2_INV_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y13__R2_INV_1 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y13__R3_BUF_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y14__R0_BUF_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R0_INV_0 (.A(tie_lo_T26Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y14__R1_BUF_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R1_INV_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R2_INV_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y14__R2_INV_1 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y14__R3_BUF_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y15__R0_BUF_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R0_INV_0 (.A(tie_lo_T26Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y15__R1_BUF_0 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R1_INV_0 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R2_INV_0 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y15__R2_INV_1 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y15__R3_BUF_0 (.A(tie_lo_T26Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y16__R0_BUF_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R0_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y16__R1_BUF_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R1_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R2_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y16__R2_INV_1 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y16__R3_BUF_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y17__R0_BUF_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R0_INV_0 (.A(tie_lo_T26Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y17__R1_BUF_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R1_INV_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R2_INV_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y17__R2_INV_1 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y17__R3_BUF_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y18__R0_BUF_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R0_INV_0 (.A(tie_lo_T26Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y18__R1_BUF_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R1_INV_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R2_INV_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y18__R2_INV_1 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y18__R3_BUF_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y19__R0_BUF_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R0_INV_0 (.A(tie_lo_T26Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y19__R1_BUF_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R1_INV_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R2_INV_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y19__R2_INV_1 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y19__R3_BUF_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y1__R0_BUF_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R0_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y1__R1_BUF_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R1_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R2_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y1__R2_INV_1 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y1__R3_BUF_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y20__R0_BUF_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R0_INV_0 (.A(tie_lo_T26Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y20__R1_BUF_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R1_INV_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R2_INV_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y20__R2_INV_1 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y20__R3_BUF_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y21__R0_BUF_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R0_INV_0 (.A(tie_lo_T26Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y21__R1_BUF_0 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R1_INV_0 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R2_INV_0 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y21__R2_INV_1 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y21__R3_BUF_0 (.A(tie_lo_T26Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y22__R0_BUF_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R0_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y22__R1_BUF_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R1_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R2_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y22__R2_INV_1 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y22__R3_BUF_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y23__R0_BUF_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R0_INV_0 (.A(tie_lo_T26Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y23__R1_BUF_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R1_INV_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R2_INV_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y23__R2_INV_1 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y23__R3_BUF_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y24__R0_BUF_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R0_INV_0 (.A(tie_lo_T26Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y24__R1_BUF_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R1_INV_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R2_INV_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y24__R2_INV_1 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y24__R3_BUF_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y25__R0_BUF_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R0_INV_0 (.A(tie_lo_T26Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y25__R1_BUF_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R1_INV_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R2_INV_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y25__R2_INV_1 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y25__R3_BUF_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y26__R0_BUF_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R0_INV_0 (.A(tie_lo_T26Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y26__R1_BUF_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R1_INV_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R2_INV_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y26__R2_INV_1 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y26__R3_BUF_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y27__R0_BUF_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R0_INV_0 (.A(tie_lo_T26Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y27__R1_BUF_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R1_INV_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R2_INV_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y27__R2_INV_1 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y27__R3_BUF_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y28__R0_BUF_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R0_INV_0 (.A(tie_lo_T26Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y28__R1_BUF_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R1_INV_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R2_INV_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y28__R2_INV_1 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y28__R3_BUF_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y29__R0_BUF_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R0_INV_0 (.A(tie_lo_T26Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y29__R1_BUF_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R1_INV_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R2_INV_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y29__R2_INV_1 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y29__R3_BUF_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y2__R0_BUF_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R0_INV_0 (.A(tie_lo_T26Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y2__R1_BUF_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R1_INV_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R2_INV_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y2__R2_INV_1 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y2__R3_BUF_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y30__R0_BUF_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R0_INV_0 (.A(tie_lo_T26Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y30__R1_BUF_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R1_INV_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R2_INV_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y30__R2_INV_1 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y30__R3_BUF_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y31__R0_BUF_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R0_INV_0 (.A(tie_lo_T26Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y31__R1_BUF_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R1_INV_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R2_INV_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y31__R2_INV_1 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y31__R3_BUF_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y32__R0_BUF_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R0_INV_0 (.A(tie_lo_T26Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y32__R1_BUF_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R1_INV_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R2_INV_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y32__R2_INV_1 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y32__R3_BUF_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y33__R0_BUF_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R0_INV_0 (.A(tie_lo_T26Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y33__R1_BUF_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R1_INV_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R2_INV_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y33__R2_INV_1 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y33__R3_BUF_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y34__R0_BUF_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R0_INV_0 (.A(tie_lo_T26Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y34__R1_BUF_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R1_INV_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R2_INV_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y34__R2_INV_1 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y34__R3_BUF_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y35__R0_BUF_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R0_INV_0 (.A(tie_lo_T26Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y35__R1_BUF_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R1_INV_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R2_INV_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y35__R2_INV_1 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y35__R3_BUF_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y36__R0_BUF_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R0_INV_0 (.A(tie_lo_T26Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y36__R1_BUF_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R1_INV_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R2_INV_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y36__R2_INV_1 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y36__R3_BUF_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y37__R0_BUF_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R0_INV_0 (.A(tie_lo_T26Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y37__R1_BUF_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R1_INV_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R2_INV_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y37__R2_INV_1 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y37__R3_BUF_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y38__R0_BUF_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R0_INV_0 (.A(tie_lo_T26Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y38__R1_BUF_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R1_INV_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R2_INV_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y38__R2_INV_1 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y38__R3_BUF_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y39__R0_BUF_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R0_INV_0 (.A(tie_lo_T26Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y39__R1_BUF_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R1_INV_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R2_INV_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y39__R2_INV_1 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y39__R3_BUF_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y3__R0_BUF_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R0_INV_0 (.A(tie_lo_T26Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y3__R1_BUF_0 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R1_INV_0 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R2_INV_0 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y3__R2_INV_1 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y3__R3_BUF_0 (.A(tie_lo_T26Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y40__R0_BUF_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R0_INV_0 (.A(tie_lo_T26Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y40__R1_BUF_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R1_INV_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R2_INV_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y40__R2_INV_1 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y40__R3_BUF_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y41__R0_BUF_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R0_INV_0 (.A(tie_lo_T26Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y41__R1_BUF_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R1_INV_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R2_INV_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y41__R2_INV_1 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y41__R3_BUF_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y42__R0_BUF_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R0_INV_0 (.A(tie_lo_T26Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y42__R1_BUF_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R1_INV_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R2_INV_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y42__R2_INV_1 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y42__R3_BUF_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y43__R0_BUF_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R0_INV_0 (.A(tie_lo_T26Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y43__R1_BUF_0 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R1_INV_0 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R2_INV_0 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y43__R2_INV_1 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y43__R3_BUF_0 (.A(tie_lo_T26Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y44__R0_BUF_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R0_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y44__R1_BUF_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R1_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R2_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y44__R2_INV_1 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y44__R3_BUF_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y45__R0_BUF_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R0_INV_0 (.A(tie_lo_T26Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y45__R1_BUF_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R1_INV_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R2_INV_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y45__R2_INV_1 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y45__R3_BUF_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y46__R0_BUF_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R0_INV_0 (.A(tie_lo_T26Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y46__R1_BUF_0 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R1_INV_0 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R2_INV_0 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y46__R2_INV_1 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y46__R3_BUF_0 (.A(tie_lo_T26Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y47__R0_BUF_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R0_INV_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y47__R1_BUF_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R1_INV_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R2_INV_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y47__R2_INV_1 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y47__R3_BUF_0 (.A(tie_lo_T26Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y48__R0_BUF_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R0_INV_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y48__R1_BUF_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R1_INV_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R2_INV_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y48__R2_INV_1 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y48__R3_BUF_0 (.A(tie_lo_T26Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y49__R0_BUF_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R0_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y49__R1_BUF_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R1_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R2_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y49__R2_INV_1 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y49__R3_BUF_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y4__R0_BUF_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R0_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y4__R1_BUF_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R1_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R2_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y4__R2_INV_1 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y4__R3_BUF_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y50__R0_BUF_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R0_INV_0 (.A(tie_lo_T26Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y50__R1_BUF_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R1_INV_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R2_INV_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y50__R2_INV_1 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y50__R3_BUF_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y51__R0_BUF_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R0_INV_0 (.A(tie_lo_T26Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y51__R1_BUF_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R1_INV_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R2_INV_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y51__R2_INV_1 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y51__R3_BUF_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y52__R0_BUF_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R0_INV_0 (.A(tie_lo_T26Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y52__R1_BUF_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R1_INV_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R2_INV_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y52__R2_INV_1 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y52__R3_BUF_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y53__R0_BUF_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R0_INV_0 (.A(tie_lo_T26Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y53__R1_BUF_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R1_INV_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R2_INV_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y53__R2_INV_1 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y53__R3_BUF_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y54__R0_BUF_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R0_INV_0 (.A(tie_lo_T26Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y54__R1_BUF_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R1_INV_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R2_INV_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y54__R2_INV_1 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y54__R3_BUF_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y55__R0_BUF_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R0_INV_0 (.A(tie_lo_T26Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y55__R1_BUF_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R1_INV_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R2_INV_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y55__R2_INV_1 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y55__R3_BUF_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y56__R0_BUF_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R0_INV_0 (.A(tie_lo_T26Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y56__R1_BUF_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R1_INV_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R2_INV_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y56__R2_INV_1 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y56__R3_BUF_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y57__R0_BUF_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R0_INV_0 (.A(tie_lo_T26Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y57__R1_BUF_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R1_INV_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R2_INV_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y57__R2_INV_1 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y57__R3_BUF_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y58__R0_BUF_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R0_INV_0 (.A(tie_lo_T26Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y58__R1_BUF_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R1_INV_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R2_INV_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y58__R2_INV_1 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y58__R3_BUF_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y59__R0_BUF_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R0_INV_0 (.A(tie_lo_T26Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y59__R1_BUF_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R1_INV_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R2_INV_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y59__R2_INV_1 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y59__R3_BUF_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y5__R0_BUF_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R0_INV_0 (.A(tie_lo_T26Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y5__R1_BUF_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R1_INV_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R2_INV_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y5__R2_INV_1 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y5__R3_BUF_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y60__R0_BUF_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R0_INV_0 (.A(tie_lo_T26Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y60__R1_BUF_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R1_INV_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R2_INV_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y60__R2_INV_1 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y60__R3_BUF_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y61__R0_BUF_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R0_INV_0 (.A(tie_lo_T26Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y61__R1_BUF_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R1_INV_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R2_INV_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y61__R2_INV_1 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y61__R3_BUF_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y62__R0_BUF_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R0_INV_0 (.A(tie_lo_T26Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y62__R1_BUF_0 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R1_INV_0 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R2_INV_0 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y62__R2_INV_1 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y62__R3_BUF_0 (.A(tie_lo_T26Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y63__R0_BUF_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R0_INV_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y63__R1_BUF_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R1_INV_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R2_INV_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y63__R2_INV_1 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y63__R3_BUF_0 (.A(tie_lo_T26Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y64__R0_BUF_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R0_INV_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y64__R1_BUF_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R1_INV_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R2_INV_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y64__R2_INV_1 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y64__R3_BUF_0 (.A(tie_lo_T26Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y65__R0_BUF_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R0_INV_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y65__R1_BUF_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R1_INV_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R2_INV_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y65__R2_INV_1 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y65__R3_BUF_0 (.A(tie_lo_T26Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y66__R0_BUF_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R0_INV_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y66__R1_BUF_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R1_INV_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R2_INV_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y66__R2_INV_1 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y66__R3_BUF_0 (.A(tie_lo_T26Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y67__R0_BUF_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R0_INV_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y67__R1_BUF_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R1_INV_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R2_INV_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y67__R2_INV_1 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y67__R3_BUF_0 (.A(tie_lo_T26Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y68__R0_BUF_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R0_INV_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y68__R1_BUF_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R1_INV_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R2_INV_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y68__R2_INV_1 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y68__R3_BUF_0 (.A(tie_lo_T26Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y69__R0_BUF_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R0_INV_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y69__R1_BUF_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R1_INV_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R2_INV_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y69__R2_INV_1 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y69__R3_BUF_0 (.A(tie_lo_T26Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y6__R0_BUF_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R0_INV_0 (.A(tie_lo_T26Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y6__R1_BUF_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R1_INV_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R2_INV_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y6__R2_INV_1 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y6__R3_BUF_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y70__R0_BUF_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R0_INV_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y70__R1_BUF_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R1_INV_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R2_INV_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y70__R2_INV_1 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y70__R3_BUF_0 (.A(tie_lo_T26Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y71__R0_BUF_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R0_INV_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y71__R1_BUF_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R1_INV_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R2_INV_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y71__R2_INV_1 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y71__R3_BUF_0 (.A(tie_lo_T26Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y72__R0_BUF_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R0_INV_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y72__R1_BUF_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R1_INV_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R2_INV_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y72__R2_INV_1 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y72__R3_BUF_0 (.A(tie_lo_T26Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y73__R0_BUF_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R0_INV_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y73__R1_BUF_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R1_INV_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R2_INV_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y73__R2_INV_1 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y73__R3_BUF_0 (.A(tie_lo_T26Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y74__R0_BUF_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R0_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y74__R1_BUF_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R1_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R2_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y74__R2_INV_1 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y74__R3_BUF_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y75__R0_BUF_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R0_INV_0 (.A(tie_lo_T26Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y75__R1_BUF_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R1_INV_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R2_INV_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y75__R2_INV_1 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y75__R3_BUF_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y76__R0_BUF_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R0_INV_0 (.A(tie_lo_T26Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y76__R1_BUF_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R1_INV_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R2_INV_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y76__R2_INV_1 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y76__R3_BUF_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y77__R0_BUF_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R0_INV_0 (.A(tie_lo_T26Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y77__R1_BUF_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R1_INV_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R2_INV_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y77__R2_INV_1 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y77__R3_BUF_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y78__R0_BUF_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R0_INV_0 (.A(tie_lo_T26Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y78__R1_BUF_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R1_INV_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R2_INV_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y78__R2_INV_1 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y78__R3_BUF_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y79__R0_BUF_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R0_INV_0 (.A(tie_lo_T26Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y79__R1_BUF_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R1_INV_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R2_INV_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y79__R2_INV_1 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y79__R3_BUF_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y7__R0_BUF_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R0_INV_0 (.A(tie_lo_T26Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y7__R1_BUF_0 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R1_INV_0 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R2_INV_0 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y7__R2_INV_1 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y7__R3_BUF_0 (.A(tie_lo_T26Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y80__R0_BUF_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R0_INV_0 (.A(tie_lo_T26Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y80__R1_BUF_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R1_INV_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R2_INV_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y80__R2_INV_1 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y80__R3_BUF_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y81__R0_BUF_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R0_INV_0 (.A(tie_lo_T26Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y81__R1_BUF_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R1_INV_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R2_INV_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y81__R2_INV_1 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y81__R3_BUF_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y82__R0_BUF_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R0_INV_0 (.A(tie_lo_T26Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y82__R1_BUF_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R1_INV_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R2_INV_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y82__R2_INV_1 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y82__R3_BUF_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y83__R0_BUF_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R0_INV_0 (.A(tie_lo_T26Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y83__R1_BUF_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R1_INV_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R2_INV_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y83__R2_INV_1 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y83__R3_BUF_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y84__R0_BUF_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R0_INV_0 (.A(tie_lo_T26Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y84__R1_BUF_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R1_INV_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R2_INV_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y84__R2_INV_1 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y84__R3_BUF_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y85__R0_BUF_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R0_INV_0 (.A(tie_lo_T26Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y85__R1_BUF_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R1_INV_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R2_INV_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y85__R2_INV_1 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y85__R3_BUF_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y86__R0_BUF_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R0_INV_0 (.A(tie_lo_T26Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y86__R1_BUF_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R1_INV_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R2_INV_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y86__R2_INV_1 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y86__R3_BUF_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y87__R0_BUF_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R0_INV_0 (.A(tie_lo_T26Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y87__R1_BUF_0 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R1_INV_0 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R2_INV_0 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y87__R2_INV_1 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y87__R3_BUF_0 (.A(tie_lo_T26Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y88__R0_BUF_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R0_INV_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y88__R1_BUF_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R1_INV_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R2_INV_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y88__R2_INV_1 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y88__R3_BUF_0 (.A(tie_lo_T26Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y89__R0_BUF_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R0_INV_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y89__R1_BUF_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R1_INV_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R2_INV_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y89__R2_INV_1 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y89__R3_BUF_0 (.A(tie_lo_T26Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y8__R0_BUF_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R0_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y8__R1_BUF_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R1_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R2_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y8__R2_INV_1 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y8__R3_BUF_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y9__R0_BUF_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R0_INV_0 (.A(tie_lo_T26Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y9__R1_BUF_0 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R1_INV_0 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T26Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R2_INV_0 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T26Y9__R2_INV_1 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T26Y9__R3_BUF_0 (.A(tie_lo_T26Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y0__R0_BUF_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R0_INV_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y0__R1_BUF_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R1_INV_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R2_INV_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y0__R2_INV_1 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y0__R3_BUF_0 (.A(tie_lo_T27Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y10__R0_BUF_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R0_INV_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y10__R1_BUF_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R1_INV_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R2_INV_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y10__R2_INV_1 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y10__R3_BUF_0 (.A(tie_lo_T27Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y11__R0_BUF_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R0_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y11__R1_BUF_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R1_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R2_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y11__R2_INV_1 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y11__R3_BUF_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y12__R0_BUF_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R0_INV_0 (.A(tie_lo_T27Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y12__R1_BUF_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R1_INV_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R2_INV_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y12__R2_INV_1 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y12__R3_BUF_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y13__R0_BUF_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R0_INV_0 (.A(tie_lo_T27Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y13__R1_BUF_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R1_INV_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R2_INV_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y13__R2_INV_1 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y13__R3_BUF_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y14__R0_BUF_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R0_INV_0 (.A(tie_lo_T27Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y14__R1_BUF_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R1_INV_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R2_INV_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y14__R2_INV_1 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y14__R3_BUF_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y15__R0_BUF_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R0_INV_0 (.A(tie_lo_T27Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y15__R1_BUF_0 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R1_INV_0 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R2_INV_0 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y15__R2_INV_1 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y15__R3_BUF_0 (.A(tie_lo_T27Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y16__R0_BUF_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R0_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y16__R1_BUF_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R1_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R2_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y16__R2_INV_1 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y16__R3_BUF_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y17__R0_BUF_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R0_INV_0 (.A(tie_lo_T27Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y17__R1_BUF_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R1_INV_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R2_INV_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y17__R2_INV_1 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y17__R3_BUF_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y18__R0_BUF_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R0_INV_0 (.A(tie_lo_T27Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y18__R1_BUF_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R1_INV_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R2_INV_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y18__R2_INV_1 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y18__R3_BUF_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y19__R0_BUF_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R0_INV_0 (.A(tie_lo_T27Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y19__R1_BUF_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R1_INV_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R2_INV_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y19__R2_INV_1 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y19__R3_BUF_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y1__R0_BUF_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R0_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y1__R1_BUF_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R1_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R2_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y1__R2_INV_1 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y1__R3_BUF_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y20__R0_BUF_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R0_INV_0 (.A(tie_lo_T27Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y20__R1_BUF_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R1_INV_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R2_INV_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y20__R2_INV_1 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y20__R3_BUF_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y21__R0_BUF_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R0_INV_0 (.A(tie_lo_T27Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y21__R1_BUF_0 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R1_INV_0 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R2_INV_0 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y21__R2_INV_1 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y21__R3_BUF_0 (.A(tie_lo_T27Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y22__R0_BUF_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R0_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y22__R1_BUF_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R1_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R2_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y22__R2_INV_1 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y22__R3_BUF_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y23__R0_BUF_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R0_INV_0 (.A(tie_lo_T27Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y23__R1_BUF_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R1_INV_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R2_INV_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y23__R2_INV_1 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y23__R3_BUF_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y24__R0_BUF_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R0_INV_0 (.A(tie_lo_T27Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y24__R1_BUF_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R1_INV_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R2_INV_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y24__R2_INV_1 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y24__R3_BUF_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y25__R0_BUF_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R0_INV_0 (.A(tie_lo_T27Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y25__R1_BUF_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R1_INV_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R2_INV_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y25__R2_INV_1 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y25__R3_BUF_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y26__R0_BUF_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R0_INV_0 (.A(tie_lo_T27Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y26__R1_BUF_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R1_INV_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R2_INV_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y26__R2_INV_1 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y26__R3_BUF_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y27__R0_BUF_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R0_INV_0 (.A(tie_lo_T27Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y27__R1_BUF_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R1_INV_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R2_INV_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y27__R2_INV_1 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y27__R3_BUF_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y28__R0_BUF_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R0_INV_0 (.A(tie_lo_T27Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y28__R1_BUF_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R1_INV_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R2_INV_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y28__R2_INV_1 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y28__R3_BUF_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y29__R0_BUF_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R0_INV_0 (.A(tie_lo_T27Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y29__R1_BUF_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R1_INV_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R2_INV_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y29__R2_INV_1 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y29__R3_BUF_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y2__R0_BUF_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R0_INV_0 (.A(tie_lo_T27Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y2__R1_BUF_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R1_INV_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R2_INV_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y2__R2_INV_1 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y2__R3_BUF_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y30__R0_BUF_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R0_INV_0 (.A(tie_lo_T27Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y30__R1_BUF_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R1_INV_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R2_INV_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y30__R2_INV_1 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y30__R3_BUF_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y31__R0_BUF_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R0_INV_0 (.A(tie_lo_T27Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y31__R1_BUF_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R1_INV_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R2_INV_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y31__R2_INV_1 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y31__R3_BUF_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y32__R0_BUF_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R0_INV_0 (.A(tie_lo_T27Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y32__R1_BUF_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R1_INV_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R2_INV_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y32__R2_INV_1 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y32__R3_BUF_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y33__R0_BUF_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R0_INV_0 (.A(tie_lo_T27Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y33__R1_BUF_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R1_INV_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R2_INV_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y33__R2_INV_1 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y33__R3_BUF_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y34__R0_BUF_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R0_INV_0 (.A(tie_lo_T27Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y34__R1_BUF_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R1_INV_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R2_INV_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y34__R2_INV_1 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y34__R3_BUF_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y35__R0_BUF_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R0_INV_0 (.A(tie_lo_T27Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y35__R1_BUF_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R1_INV_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R2_INV_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y35__R2_INV_1 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y35__R3_BUF_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y36__R0_BUF_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R0_INV_0 (.A(tie_lo_T27Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y36__R1_BUF_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R1_INV_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R2_INV_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y36__R2_INV_1 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y36__R3_BUF_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y37__R0_BUF_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R0_INV_0 (.A(tie_lo_T27Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y37__R1_BUF_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R1_INV_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R2_INV_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y37__R2_INV_1 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y37__R3_BUF_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y38__R0_BUF_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R0_INV_0 (.A(tie_lo_T27Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y38__R1_BUF_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R1_INV_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R2_INV_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y38__R2_INV_1 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y38__R3_BUF_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y39__R0_BUF_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R0_INV_0 (.A(tie_lo_T27Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y39__R1_BUF_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R1_INV_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R2_INV_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y39__R2_INV_1 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y39__R3_BUF_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y3__R0_BUF_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R0_INV_0 (.A(tie_lo_T27Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y3__R1_BUF_0 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R1_INV_0 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R2_INV_0 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y3__R2_INV_1 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y3__R3_BUF_0 (.A(tie_lo_T27Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y40__R0_BUF_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R0_INV_0 (.A(tie_lo_T27Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y40__R1_BUF_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R1_INV_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R2_INV_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y40__R2_INV_1 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y40__R3_BUF_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y41__R0_BUF_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R0_INV_0 (.A(tie_lo_T27Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y41__R1_BUF_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R1_INV_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R2_INV_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y41__R2_INV_1 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y41__R3_BUF_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y42__R0_BUF_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R0_INV_0 (.A(tie_lo_T27Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y42__R1_BUF_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R1_INV_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R2_INV_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y42__R2_INV_1 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y42__R3_BUF_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y43__R0_BUF_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R0_INV_0 (.A(tie_lo_T27Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y43__R1_BUF_0 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R1_INV_0 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R2_INV_0 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y43__R2_INV_1 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y43__R3_BUF_0 (.A(tie_lo_T27Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y44__R0_BUF_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R0_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y44__R1_BUF_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R1_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R2_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y44__R2_INV_1 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y44__R3_BUF_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y45__R0_BUF_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R0_INV_0 (.A(tie_lo_T27Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y45__R1_BUF_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R1_INV_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R2_INV_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y45__R2_INV_1 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y45__R3_BUF_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y46__R0_BUF_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R0_INV_0 (.A(tie_lo_T27Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y46__R1_BUF_0 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R1_INV_0 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R2_INV_0 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y46__R2_INV_1 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y46__R3_BUF_0 (.A(tie_lo_T27Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y47__R0_BUF_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R0_INV_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y47__R1_BUF_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R1_INV_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R2_INV_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y47__R2_INV_1 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y47__R3_BUF_0 (.A(tie_lo_T27Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y48__R0_BUF_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R0_INV_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y48__R1_BUF_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R1_INV_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R2_INV_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y48__R2_INV_1 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y48__R3_BUF_0 (.A(tie_lo_T27Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y49__R0_BUF_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R0_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y49__R1_BUF_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R1_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R2_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y49__R2_INV_1 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y49__R3_BUF_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y4__R0_BUF_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R0_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y4__R1_BUF_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R1_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R2_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y4__R2_INV_1 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y4__R3_BUF_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y50__R0_BUF_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R0_INV_0 (.A(tie_lo_T27Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y50__R1_BUF_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R1_INV_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R2_INV_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y50__R2_INV_1 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y50__R3_BUF_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y51__R0_BUF_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R0_INV_0 (.A(tie_lo_T27Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y51__R1_BUF_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R1_INV_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R2_INV_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y51__R2_INV_1 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y51__R3_BUF_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y52__R0_BUF_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R0_INV_0 (.A(tie_lo_T27Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y52__R1_BUF_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R1_INV_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R2_INV_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y52__R2_INV_1 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y52__R3_BUF_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y53__R0_BUF_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R0_INV_0 (.A(tie_lo_T27Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y53__R1_BUF_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R1_INV_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R2_INV_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y53__R2_INV_1 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y53__R3_BUF_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y54__R0_BUF_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R0_INV_0 (.A(tie_lo_T27Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y54__R1_BUF_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R1_INV_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R2_INV_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y54__R2_INV_1 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y54__R3_BUF_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y55__R0_BUF_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R0_INV_0 (.A(tie_lo_T27Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y55__R1_BUF_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R1_INV_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R2_INV_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y55__R2_INV_1 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y55__R3_BUF_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y56__R0_BUF_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R0_INV_0 (.A(tie_lo_T27Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y56__R1_BUF_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R1_INV_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R2_INV_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y56__R2_INV_1 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y56__R3_BUF_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y57__R0_BUF_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R0_INV_0 (.A(tie_lo_T27Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y57__R1_BUF_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R1_INV_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R2_INV_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y57__R2_INV_1 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y57__R3_BUF_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y58__R0_BUF_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R0_INV_0 (.A(tie_lo_T27Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y58__R1_BUF_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R1_INV_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R2_INV_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y58__R2_INV_1 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y58__R3_BUF_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y59__R0_BUF_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R0_INV_0 (.A(tie_lo_T27Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y59__R1_BUF_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R1_INV_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R2_INV_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y59__R2_INV_1 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y59__R3_BUF_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y5__R0_BUF_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R0_INV_0 (.A(tie_lo_T27Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y5__R1_BUF_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R1_INV_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R2_INV_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y5__R2_INV_1 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y5__R3_BUF_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y60__R0_BUF_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R0_INV_0 (.A(tie_lo_T27Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y60__R1_BUF_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R1_INV_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R2_INV_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y60__R2_INV_1 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y60__R3_BUF_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y61__R0_BUF_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R0_INV_0 (.A(tie_lo_T27Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y61__R1_BUF_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R1_INV_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R2_INV_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y61__R2_INV_1 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y61__R3_BUF_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y62__R0_BUF_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R0_INV_0 (.A(tie_lo_T27Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y62__R1_BUF_0 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R1_INV_0 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R2_INV_0 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y62__R2_INV_1 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y62__R3_BUF_0 (.A(tie_lo_T27Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y63__R0_BUF_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R0_INV_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y63__R1_BUF_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R1_INV_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R2_INV_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y63__R2_INV_1 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y63__R3_BUF_0 (.A(tie_lo_T27Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y64__R0_BUF_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R0_INV_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y64__R1_BUF_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R1_INV_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R2_INV_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y64__R2_INV_1 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y64__R3_BUF_0 (.A(tie_lo_T27Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y65__R0_BUF_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R0_INV_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y65__R1_BUF_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R1_INV_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R2_INV_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y65__R2_INV_1 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y65__R3_BUF_0 (.A(tie_lo_T27Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y66__R0_BUF_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R0_INV_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y66__R1_BUF_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R1_INV_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R2_INV_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y66__R2_INV_1 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y66__R3_BUF_0 (.A(tie_lo_T27Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y67__R0_BUF_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R0_INV_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y67__R1_BUF_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R1_INV_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R2_INV_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y67__R2_INV_1 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y67__R3_BUF_0 (.A(tie_lo_T27Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y68__R0_BUF_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R0_INV_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y68__R1_BUF_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R1_INV_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R2_INV_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y68__R2_INV_1 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y68__R3_BUF_0 (.A(tie_lo_T27Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y69__R0_BUF_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R0_INV_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y69__R1_BUF_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R1_INV_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R2_INV_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y69__R2_INV_1 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y69__R3_BUF_0 (.A(tie_lo_T27Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y6__R0_BUF_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R0_INV_0 (.A(tie_lo_T27Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y6__R1_BUF_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R1_INV_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R2_INV_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y6__R2_INV_1 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y6__R3_BUF_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y70__R0_BUF_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R0_INV_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y70__R1_BUF_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R1_INV_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R2_INV_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y70__R2_INV_1 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y70__R3_BUF_0 (.A(tie_lo_T27Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y71__R0_BUF_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R0_INV_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y71__R1_BUF_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R1_INV_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R2_INV_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y71__R2_INV_1 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y71__R3_BUF_0 (.A(tie_lo_T27Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y72__R0_BUF_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R0_INV_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y72__R1_BUF_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R1_INV_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R2_INV_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y72__R2_INV_1 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y72__R3_BUF_0 (.A(tie_lo_T27Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y73__R0_BUF_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R0_INV_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y73__R1_BUF_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R1_INV_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R2_INV_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y73__R2_INV_1 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y73__R3_BUF_0 (.A(tie_lo_T27Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y74__R0_BUF_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R0_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y74__R1_BUF_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R1_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R2_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y74__R2_INV_1 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y74__R3_BUF_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y75__R0_BUF_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R0_INV_0 (.A(tie_lo_T27Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y75__R1_BUF_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R1_INV_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R2_INV_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y75__R2_INV_1 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y75__R3_BUF_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y76__R0_BUF_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R0_INV_0 (.A(tie_lo_T27Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y76__R1_BUF_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R1_INV_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R2_INV_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y76__R2_INV_1 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y76__R3_BUF_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y77__R0_BUF_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R0_INV_0 (.A(tie_lo_T27Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y77__R1_BUF_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R1_INV_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R2_INV_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y77__R2_INV_1 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y77__R3_BUF_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y78__R0_BUF_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R0_INV_0 (.A(tie_lo_T27Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y78__R1_BUF_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R1_INV_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R2_INV_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y78__R2_INV_1 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y78__R3_BUF_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y79__R0_BUF_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R0_INV_0 (.A(tie_lo_T27Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y79__R1_BUF_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R1_INV_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R2_INV_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y79__R2_INV_1 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y79__R3_BUF_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y7__R0_BUF_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R0_INV_0 (.A(tie_lo_T27Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y7__R1_BUF_0 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R1_INV_0 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R2_INV_0 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y7__R2_INV_1 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y7__R3_BUF_0 (.A(tie_lo_T27Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y80__R0_BUF_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R0_INV_0 (.A(tie_lo_T27Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y80__R1_BUF_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R1_INV_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R2_INV_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y80__R2_INV_1 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y80__R3_BUF_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y81__R0_BUF_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R0_INV_0 (.A(tie_lo_T27Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y81__R1_BUF_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R1_INV_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R2_INV_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y81__R2_INV_1 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y81__R3_BUF_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y82__R0_BUF_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R0_INV_0 (.A(tie_lo_T27Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y82__R1_BUF_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R1_INV_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R2_INV_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y82__R2_INV_1 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y82__R3_BUF_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y83__R0_BUF_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R0_INV_0 (.A(tie_lo_T27Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y83__R1_BUF_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R1_INV_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R2_INV_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y83__R2_INV_1 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y83__R3_BUF_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y84__R0_BUF_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R0_INV_0 (.A(tie_lo_T27Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y84__R1_BUF_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R1_INV_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R2_INV_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y84__R2_INV_1 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y84__R3_BUF_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y85__R0_BUF_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R0_INV_0 (.A(tie_lo_T27Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y85__R1_BUF_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R1_INV_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R2_INV_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y85__R2_INV_1 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y85__R3_BUF_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y86__R0_BUF_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R0_INV_0 (.A(tie_lo_T27Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y86__R1_BUF_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R1_INV_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R2_INV_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y86__R2_INV_1 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y86__R3_BUF_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y87__R0_BUF_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R0_INV_0 (.A(tie_lo_T27Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y87__R1_BUF_0 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R1_INV_0 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R2_INV_0 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y87__R2_INV_1 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y87__R3_BUF_0 (.A(tie_lo_T27Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y88__R0_BUF_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R0_INV_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y88__R1_BUF_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R1_INV_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R2_INV_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y88__R2_INV_1 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y88__R3_BUF_0 (.A(tie_lo_T27Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y89__R0_BUF_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R0_INV_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y89__R1_BUF_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R1_INV_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R2_INV_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y89__R2_INV_1 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y89__R3_BUF_0 (.A(tie_lo_T27Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y8__R0_BUF_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R0_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y8__R1_BUF_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R1_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R2_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y8__R2_INV_1 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y8__R3_BUF_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y9__R0_BUF_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R0_INV_0 (.A(tie_lo_T27Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y9__R1_BUF_0 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R1_INV_0 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T27Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R2_INV_0 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T27Y9__R2_INV_1 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T27Y9__R3_BUF_0 (.A(tie_lo_T27Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y0__R0_BUF_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R0_INV_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y0__R1_BUF_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R1_INV_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R2_INV_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y0__R2_INV_1 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y0__R3_BUF_0 (.A(tie_lo_T28Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y10__R0_BUF_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R0_INV_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y10__R1_BUF_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R1_INV_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R2_INV_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y10__R2_INV_1 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y10__R3_BUF_0 (.A(tie_lo_T28Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y11__R0_BUF_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R0_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y11__R1_BUF_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R1_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R2_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y11__R2_INV_1 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y11__R3_BUF_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y12__R0_BUF_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R0_INV_0 (.A(tie_lo_T28Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y12__R1_BUF_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R1_INV_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R2_INV_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y12__R2_INV_1 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y12__R3_BUF_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y13__R0_BUF_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R0_INV_0 (.A(tie_lo_T28Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y13__R1_BUF_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R1_INV_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R2_INV_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y13__R2_INV_1 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y13__R3_BUF_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y14__R0_BUF_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R0_INV_0 (.A(tie_lo_T28Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y14__R1_BUF_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R1_INV_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R2_INV_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y14__R2_INV_1 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y14__R3_BUF_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y15__R0_BUF_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R0_INV_0 (.A(tie_lo_T28Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y15__R1_BUF_0 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R1_INV_0 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R2_INV_0 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y15__R2_INV_1 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y15__R3_BUF_0 (.A(tie_lo_T28Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y16__R0_BUF_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R0_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y16__R1_BUF_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R1_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R2_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y16__R2_INV_1 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y16__R3_BUF_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y17__R0_BUF_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R0_INV_0 (.A(tie_lo_T28Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y17__R1_BUF_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R1_INV_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R2_INV_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y17__R2_INV_1 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y17__R3_BUF_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y18__R0_BUF_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R0_INV_0 (.A(tie_lo_T28Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y18__R1_BUF_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R1_INV_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R2_INV_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y18__R2_INV_1 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y18__R3_BUF_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y19__R0_BUF_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R0_INV_0 (.A(tie_lo_T28Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y19__R1_BUF_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R1_INV_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R2_INV_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y19__R2_INV_1 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y19__R3_BUF_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y1__R0_BUF_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R0_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y1__R1_BUF_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R1_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R2_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y1__R2_INV_1 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y1__R3_BUF_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y20__R0_BUF_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R0_INV_0 (.A(tie_lo_T28Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y20__R1_BUF_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R1_INV_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R2_INV_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y20__R2_INV_1 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y20__R3_BUF_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y21__R0_BUF_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R0_INV_0 (.A(tie_lo_T28Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y21__R1_BUF_0 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R1_INV_0 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R2_INV_0 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y21__R2_INV_1 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y21__R3_BUF_0 (.A(tie_lo_T28Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y22__R0_BUF_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R0_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y22__R1_BUF_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R1_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R2_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y22__R2_INV_1 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y22__R3_BUF_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y23__R0_BUF_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R0_INV_0 (.A(tie_lo_T28Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y23__R1_BUF_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R1_INV_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R2_INV_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y23__R2_INV_1 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y23__R3_BUF_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y24__R0_BUF_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R0_INV_0 (.A(tie_lo_T28Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y24__R1_BUF_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R1_INV_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R2_INV_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y24__R2_INV_1 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y24__R3_BUF_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y25__R0_BUF_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R0_INV_0 (.A(tie_lo_T28Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y25__R1_BUF_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R1_INV_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R2_INV_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y25__R2_INV_1 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y25__R3_BUF_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y26__R0_BUF_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R0_INV_0 (.A(tie_lo_T28Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y26__R1_BUF_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R1_INV_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R2_INV_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y26__R2_INV_1 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y26__R3_BUF_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y27__R0_BUF_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R0_INV_0 (.A(tie_lo_T28Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y27__R1_BUF_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R1_INV_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R2_INV_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y27__R2_INV_1 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y27__R3_BUF_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y28__R0_BUF_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R0_INV_0 (.A(tie_lo_T28Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y28__R1_BUF_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R1_INV_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R2_INV_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y28__R2_INV_1 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y28__R3_BUF_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y29__R0_BUF_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R0_INV_0 (.A(tie_lo_T28Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y29__R1_BUF_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R1_INV_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R2_INV_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y29__R2_INV_1 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y29__R3_BUF_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y2__R0_BUF_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R0_INV_0 (.A(tie_lo_T28Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y2__R1_BUF_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R1_INV_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R2_INV_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y2__R2_INV_1 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y2__R3_BUF_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y30__R0_BUF_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R0_INV_0 (.A(tie_lo_T28Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y30__R1_BUF_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R1_INV_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R2_INV_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y30__R2_INV_1 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y30__R3_BUF_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y31__R0_BUF_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R0_INV_0 (.A(tie_lo_T28Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y31__R1_BUF_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R1_INV_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R2_INV_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y31__R2_INV_1 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y31__R3_BUF_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y32__R0_BUF_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R0_INV_0 (.A(tie_lo_T28Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y32__R1_BUF_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R1_INV_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R2_INV_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y32__R2_INV_1 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y32__R3_BUF_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y33__R0_BUF_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R0_INV_0 (.A(tie_lo_T28Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y33__R1_BUF_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R1_INV_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R2_INV_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y33__R2_INV_1 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y33__R3_BUF_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y34__R0_BUF_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R0_INV_0 (.A(tie_lo_T28Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y34__R1_BUF_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R1_INV_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R2_INV_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y34__R2_INV_1 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y34__R3_BUF_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y35__R0_BUF_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R0_INV_0 (.A(tie_lo_T28Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y35__R1_BUF_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R1_INV_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R2_INV_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y35__R2_INV_1 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y35__R3_BUF_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y36__R0_BUF_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R0_INV_0 (.A(tie_lo_T28Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y36__R1_BUF_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R1_INV_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R2_INV_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y36__R2_INV_1 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y36__R3_BUF_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y37__R0_BUF_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R0_INV_0 (.A(tie_lo_T28Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y37__R1_BUF_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R1_INV_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R2_INV_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y37__R2_INV_1 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y37__R3_BUF_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y38__R0_BUF_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R0_INV_0 (.A(tie_lo_T28Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y38__R1_BUF_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R1_INV_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R2_INV_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y38__R2_INV_1 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y38__R3_BUF_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y39__R0_BUF_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R0_INV_0 (.A(tie_lo_T28Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y39__R1_BUF_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R1_INV_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R2_INV_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y39__R2_INV_1 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y39__R3_BUF_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y3__R0_BUF_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R0_INV_0 (.A(tie_lo_T28Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y3__R1_BUF_0 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R1_INV_0 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R2_INV_0 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y3__R2_INV_1 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y3__R3_BUF_0 (.A(tie_lo_T28Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y40__R0_BUF_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R0_INV_0 (.A(tie_lo_T28Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y40__R1_BUF_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R1_INV_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R2_INV_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y40__R2_INV_1 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y40__R3_BUF_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y41__R0_BUF_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R0_INV_0 (.A(tie_lo_T28Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y41__R1_BUF_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R1_INV_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R2_INV_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y41__R2_INV_1 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y41__R3_BUF_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y42__R0_BUF_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R0_INV_0 (.A(tie_lo_T28Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y42__R1_BUF_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R1_INV_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R2_INV_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y42__R2_INV_1 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y42__R3_BUF_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y43__R0_BUF_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R0_INV_0 (.A(tie_lo_T28Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y43__R1_BUF_0 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R1_INV_0 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R2_INV_0 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y43__R2_INV_1 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y43__R3_BUF_0 (.A(tie_lo_T28Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y44__R0_BUF_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R0_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y44__R1_BUF_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R1_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R2_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y44__R2_INV_1 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y44__R3_BUF_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y45__R0_BUF_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R0_INV_0 (.A(tie_lo_T28Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y45__R1_BUF_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R1_INV_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R2_INV_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y45__R2_INV_1 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y45__R3_BUF_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y46__R0_BUF_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R0_INV_0 (.A(tie_lo_T28Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y46__R1_BUF_0 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R1_INV_0 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R2_INV_0 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y46__R2_INV_1 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y46__R3_BUF_0 (.A(tie_lo_T28Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y47__R0_BUF_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R0_INV_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y47__R1_BUF_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R1_INV_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R2_INV_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y47__R2_INV_1 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y47__R3_BUF_0 (.A(tie_lo_T28Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y48__R0_BUF_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R0_INV_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y48__R1_BUF_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R1_INV_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R2_INV_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y48__R2_INV_1 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y48__R3_BUF_0 (.A(tie_lo_T28Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y49__R0_BUF_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R0_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y49__R1_BUF_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R1_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R2_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y49__R2_INV_1 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y49__R3_BUF_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y4__R0_BUF_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R0_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y4__R1_BUF_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R1_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R2_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y4__R2_INV_1 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y4__R3_BUF_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y50__R0_BUF_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R0_INV_0 (.A(tie_lo_T28Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y50__R1_BUF_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R1_INV_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R2_INV_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y50__R2_INV_1 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y50__R3_BUF_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y51__R0_BUF_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R0_INV_0 (.A(tie_lo_T28Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y51__R1_BUF_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R1_INV_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R2_INV_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y51__R2_INV_1 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y51__R3_BUF_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y52__R0_BUF_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R0_INV_0 (.A(tie_lo_T28Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y52__R1_BUF_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R1_INV_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R2_INV_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y52__R2_INV_1 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y52__R3_BUF_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y53__R0_BUF_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R0_INV_0 (.A(tie_lo_T28Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y53__R1_BUF_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R1_INV_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R2_INV_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y53__R2_INV_1 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y53__R3_BUF_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y54__R0_BUF_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R0_INV_0 (.A(tie_lo_T28Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y54__R1_BUF_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R1_INV_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R2_INV_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y54__R2_INV_1 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y54__R3_BUF_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y55__R0_BUF_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R0_INV_0 (.A(tie_lo_T28Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y55__R1_BUF_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R1_INV_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R2_INV_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y55__R2_INV_1 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y55__R3_BUF_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y56__R0_BUF_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R0_INV_0 (.A(tie_lo_T28Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y56__R1_BUF_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R1_INV_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R2_INV_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y56__R2_INV_1 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y56__R3_BUF_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y57__R0_BUF_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R0_INV_0 (.A(tie_lo_T28Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y57__R1_BUF_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R1_INV_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R2_INV_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y57__R2_INV_1 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y57__R3_BUF_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y58__R0_BUF_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R0_INV_0 (.A(tie_lo_T28Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y58__R1_BUF_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R1_INV_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R2_INV_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y58__R2_INV_1 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y58__R3_BUF_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y59__R0_BUF_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R0_INV_0 (.A(tie_lo_T28Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y59__R1_BUF_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R1_INV_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R2_INV_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y59__R2_INV_1 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y59__R3_BUF_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y5__R0_BUF_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R0_INV_0 (.A(tie_lo_T28Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y5__R1_BUF_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R1_INV_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R2_INV_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y5__R2_INV_1 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y5__R3_BUF_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y60__R0_BUF_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R0_INV_0 (.A(tie_lo_T28Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y60__R1_BUF_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R1_INV_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R2_INV_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y60__R2_INV_1 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y60__R3_BUF_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y61__R0_BUF_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R0_INV_0 (.A(tie_lo_T28Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y61__R1_BUF_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R1_INV_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R2_INV_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y61__R2_INV_1 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y61__R3_BUF_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y62__R0_BUF_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R0_INV_0 (.A(tie_lo_T28Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y62__R1_BUF_0 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R1_INV_0 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R2_INV_0 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y62__R2_INV_1 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y62__R3_BUF_0 (.A(tie_lo_T28Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y63__R0_BUF_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R0_INV_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y63__R1_BUF_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R1_INV_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R2_INV_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y63__R2_INV_1 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y63__R3_BUF_0 (.A(tie_lo_T28Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y64__R0_BUF_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R0_INV_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y64__R1_BUF_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R1_INV_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R2_INV_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y64__R2_INV_1 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y64__R3_BUF_0 (.A(tie_lo_T28Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y65__R0_BUF_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R0_INV_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y65__R1_BUF_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R1_INV_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R2_INV_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y65__R2_INV_1 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y65__R3_BUF_0 (.A(tie_lo_T28Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y66__R0_BUF_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R0_INV_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y66__R1_BUF_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R1_INV_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R2_INV_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y66__R2_INV_1 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y66__R3_BUF_0 (.A(tie_lo_T28Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y67__R0_BUF_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R0_INV_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y67__R1_BUF_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R1_INV_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R2_INV_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y67__R2_INV_1 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y67__R3_BUF_0 (.A(tie_lo_T28Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y68__R0_BUF_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R0_INV_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y68__R1_BUF_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R1_INV_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R2_INV_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y68__R2_INV_1 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y68__R3_BUF_0 (.A(tie_lo_T28Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y69__R0_BUF_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R0_INV_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y69__R1_BUF_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R1_INV_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R2_INV_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y69__R2_INV_1 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y69__R3_BUF_0 (.A(tie_lo_T28Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y6__R0_BUF_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R0_INV_0 (.A(tie_lo_T28Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y6__R1_BUF_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R1_INV_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R2_INV_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y6__R2_INV_1 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y6__R3_BUF_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y70__R0_BUF_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R0_INV_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y70__R1_BUF_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R1_INV_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R2_INV_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y70__R2_INV_1 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y70__R3_BUF_0 (.A(tie_lo_T28Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y71__R0_BUF_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R0_INV_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y71__R1_BUF_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R1_INV_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R2_INV_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y71__R2_INV_1 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y71__R3_BUF_0 (.A(tie_lo_T28Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y72__R0_BUF_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R0_INV_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y72__R1_BUF_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R1_INV_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R2_INV_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y72__R2_INV_1 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y72__R3_BUF_0 (.A(tie_lo_T28Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y73__R0_BUF_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R0_INV_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y73__R1_BUF_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R1_INV_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R2_INV_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y73__R2_INV_1 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y73__R3_BUF_0 (.A(tie_lo_T28Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y74__R0_BUF_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R0_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y74__R1_BUF_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R1_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R2_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y74__R2_INV_1 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y74__R3_BUF_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y75__R0_BUF_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R0_INV_0 (.A(tie_lo_T28Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y75__R1_BUF_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R1_INV_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R2_INV_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y75__R2_INV_1 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y75__R3_BUF_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y76__R0_BUF_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R0_INV_0 (.A(tie_lo_T28Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y76__R1_BUF_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R1_INV_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R2_INV_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y76__R2_INV_1 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y76__R3_BUF_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y77__R0_BUF_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R0_INV_0 (.A(tie_lo_T28Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y77__R1_BUF_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R1_INV_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R2_INV_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y77__R2_INV_1 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y77__R3_BUF_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y78__R0_BUF_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R0_INV_0 (.A(tie_lo_T28Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y78__R1_BUF_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R1_INV_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R2_INV_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y78__R2_INV_1 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y78__R3_BUF_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y79__R0_BUF_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R0_INV_0 (.A(tie_lo_T28Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y79__R1_BUF_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R1_INV_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R2_INV_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y79__R2_INV_1 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y79__R3_BUF_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y7__R0_BUF_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R0_INV_0 (.A(tie_lo_T28Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y7__R1_BUF_0 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R1_INV_0 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R2_INV_0 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y7__R2_INV_1 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y7__R3_BUF_0 (.A(tie_lo_T28Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y80__R0_BUF_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R0_INV_0 (.A(tie_lo_T28Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y80__R1_BUF_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R1_INV_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R2_INV_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y80__R2_INV_1 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y80__R3_BUF_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y81__R0_BUF_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R0_INV_0 (.A(tie_lo_T28Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y81__R1_BUF_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R1_INV_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R2_INV_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y81__R2_INV_1 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y81__R3_BUF_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y82__R0_BUF_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R0_INV_0 (.A(tie_lo_T28Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y82__R1_BUF_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R1_INV_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R2_INV_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y82__R2_INV_1 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y82__R3_BUF_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y83__R0_BUF_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R0_INV_0 (.A(tie_lo_T28Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y83__R1_BUF_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R1_INV_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R2_INV_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y83__R2_INV_1 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y83__R3_BUF_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y84__R0_BUF_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R0_INV_0 (.A(tie_lo_T28Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y84__R1_BUF_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R1_INV_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R2_INV_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y84__R2_INV_1 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y84__R3_BUF_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y85__R0_BUF_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R0_INV_0 (.A(tie_lo_T28Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y85__R1_BUF_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R1_INV_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R2_INV_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y85__R2_INV_1 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y85__R3_BUF_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y86__R0_BUF_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R0_INV_0 (.A(tie_lo_T28Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y86__R1_BUF_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R1_INV_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R2_INV_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y86__R2_INV_1 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y86__R3_BUF_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y87__R0_BUF_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R0_INV_0 (.A(tie_lo_T28Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y87__R1_BUF_0 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R1_INV_0 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R2_INV_0 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y87__R2_INV_1 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y87__R3_BUF_0 (.A(tie_lo_T28Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y88__R0_BUF_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R0_INV_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y88__R1_BUF_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R1_INV_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R2_INV_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y88__R2_INV_1 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y88__R3_BUF_0 (.A(tie_lo_T28Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y89__R0_BUF_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R0_INV_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y89__R1_BUF_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R1_INV_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R2_INV_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y89__R2_INV_1 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y89__R3_BUF_0 (.A(tie_lo_T28Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y8__R0_BUF_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R0_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y8__R1_BUF_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R1_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R2_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y8__R2_INV_1 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y8__R3_BUF_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y9__R0_BUF_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R0_INV_0 (.A(tie_lo_T28Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y9__R1_BUF_0 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R1_INV_0 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T28Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R2_INV_0 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T28Y9__R2_INV_1 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T28Y9__R3_BUF_0 (.A(tie_lo_T28Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y0__R0_BUF_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R0_INV_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y0__R1_BUF_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R1_INV_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R2_INV_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y0__R2_INV_1 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y0__R3_BUF_0 (.A(tie_lo_T29Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y10__R0_BUF_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R0_INV_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y10__R1_BUF_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R1_INV_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R2_INV_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y10__R2_INV_1 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y10__R3_BUF_0 (.A(tie_lo_T29Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y11__R0_BUF_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R0_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y11__R1_BUF_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R1_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R2_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y11__R2_INV_1 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y11__R3_BUF_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y12__R0_BUF_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R0_INV_0 (.A(tie_lo_T29Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y12__R1_BUF_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R1_INV_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R2_INV_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y12__R2_INV_1 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y12__R3_BUF_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y13__R0_BUF_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R0_INV_0 (.A(tie_lo_T29Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y13__R1_BUF_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R1_INV_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R2_INV_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y13__R2_INV_1 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y13__R3_BUF_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y14__R0_BUF_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R0_INV_0 (.A(tie_lo_T29Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y14__R1_BUF_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R1_INV_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R2_INV_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y14__R2_INV_1 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y14__R3_BUF_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y15__R0_BUF_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R0_INV_0 (.A(tie_lo_T29Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y15__R1_BUF_0 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R1_INV_0 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R2_INV_0 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y15__R2_INV_1 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y15__R3_BUF_0 (.A(tie_lo_T29Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y16__R0_BUF_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R0_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y16__R1_BUF_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R1_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R2_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y16__R2_INV_1 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y16__R3_BUF_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y17__R0_BUF_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R0_INV_0 (.A(tie_lo_T29Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y17__R1_BUF_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R1_INV_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R2_INV_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y17__R2_INV_1 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y17__R3_BUF_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y18__R0_BUF_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R0_INV_0 (.A(tie_lo_T29Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y18__R1_BUF_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R1_INV_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R2_INV_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y18__R2_INV_1 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y18__R3_BUF_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y19__R0_BUF_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R0_INV_0 (.A(tie_lo_T29Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y19__R1_BUF_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R1_INV_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R2_INV_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y19__R2_INV_1 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y19__R3_BUF_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y1__R0_BUF_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R0_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y1__R1_BUF_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R1_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R2_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y1__R2_INV_1 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y1__R3_BUF_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y20__R0_BUF_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R0_INV_0 (.A(tie_lo_T29Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y20__R1_BUF_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R1_INV_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R2_INV_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y20__R2_INV_1 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y20__R3_BUF_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y21__R0_BUF_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R0_INV_0 (.A(tie_lo_T29Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y21__R1_BUF_0 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R1_INV_0 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R2_INV_0 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y21__R2_INV_1 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y21__R3_BUF_0 (.A(tie_lo_T29Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y22__R0_BUF_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R0_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y22__R1_BUF_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R1_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R2_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y22__R2_INV_1 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y22__R3_BUF_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y23__R0_BUF_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R0_INV_0 (.A(tie_lo_T29Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y23__R1_BUF_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R1_INV_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R2_INV_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y23__R2_INV_1 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y23__R3_BUF_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y24__R0_BUF_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R0_INV_0 (.A(tie_lo_T29Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y24__R1_BUF_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R1_INV_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R2_INV_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y24__R2_INV_1 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y24__R3_BUF_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y25__R0_BUF_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R0_INV_0 (.A(tie_lo_T29Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y25__R1_BUF_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R1_INV_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R2_INV_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y25__R2_INV_1 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y25__R3_BUF_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y26__R0_BUF_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R0_INV_0 (.A(tie_lo_T29Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y26__R1_BUF_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R1_INV_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R2_INV_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y26__R2_INV_1 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y26__R3_BUF_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y27__R0_BUF_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R0_INV_0 (.A(tie_lo_T29Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y27__R1_BUF_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R1_INV_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R2_INV_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y27__R2_INV_1 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y27__R3_BUF_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y28__R0_BUF_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R0_INV_0 (.A(tie_lo_T29Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y28__R1_BUF_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R1_INV_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R2_INV_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y28__R2_INV_1 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y28__R3_BUF_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y29__R0_BUF_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R0_INV_0 (.A(tie_lo_T29Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y29__R1_BUF_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R1_INV_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R2_INV_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y29__R2_INV_1 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y29__R3_BUF_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y2__R0_BUF_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R0_INV_0 (.A(tie_lo_T29Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y2__R1_BUF_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R1_INV_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R2_INV_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y2__R2_INV_1 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y2__R3_BUF_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y30__R0_BUF_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R0_INV_0 (.A(tie_lo_T29Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y30__R1_BUF_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R1_INV_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R2_INV_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y30__R2_INV_1 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y30__R3_BUF_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y31__R0_BUF_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R0_INV_0 (.A(tie_lo_T29Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y31__R1_BUF_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R1_INV_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R2_INV_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y31__R2_INV_1 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y31__R3_BUF_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y32__R0_BUF_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R0_INV_0 (.A(tie_lo_T29Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y32__R1_BUF_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R1_INV_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R2_INV_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y32__R2_INV_1 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y32__R3_BUF_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y33__R0_BUF_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R0_INV_0 (.A(tie_lo_T29Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y33__R1_BUF_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R1_INV_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R2_INV_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y33__R2_INV_1 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y33__R3_BUF_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y34__R0_BUF_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R0_INV_0 (.A(tie_lo_T29Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y34__R1_BUF_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R1_INV_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R2_INV_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y34__R2_INV_1 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y34__R3_BUF_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y35__R0_BUF_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R0_INV_0 (.A(tie_lo_T29Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y35__R1_BUF_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R1_INV_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R2_INV_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y35__R2_INV_1 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y35__R3_BUF_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y36__R0_BUF_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R0_INV_0 (.A(tie_lo_T29Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y36__R1_BUF_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R1_INV_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R2_INV_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y36__R2_INV_1 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y36__R3_BUF_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y37__R0_BUF_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R0_INV_0 (.A(tie_lo_T29Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y37__R1_BUF_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R1_INV_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R2_INV_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y37__R2_INV_1 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y37__R3_BUF_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y38__R0_BUF_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R0_INV_0 (.A(tie_lo_T29Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y38__R1_BUF_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R1_INV_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R2_INV_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y38__R2_INV_1 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y38__R3_BUF_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y39__R0_BUF_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R0_INV_0 (.A(tie_lo_T29Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y39__R1_BUF_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R1_INV_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R2_INV_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y39__R2_INV_1 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y39__R3_BUF_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y3__R0_BUF_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R0_INV_0 (.A(tie_lo_T29Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y3__R1_BUF_0 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R1_INV_0 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R2_INV_0 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y3__R2_INV_1 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y3__R3_BUF_0 (.A(tie_lo_T29Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y40__R0_BUF_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R0_INV_0 (.A(tie_lo_T29Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y40__R1_BUF_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R1_INV_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R2_INV_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y40__R2_INV_1 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y40__R3_BUF_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y41__R0_BUF_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R0_INV_0 (.A(tie_lo_T29Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y41__R1_BUF_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R1_INV_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R2_INV_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y41__R2_INV_1 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y41__R3_BUF_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y42__R0_BUF_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R0_INV_0 (.A(tie_lo_T29Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y42__R1_BUF_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R1_INV_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R2_INV_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y42__R2_INV_1 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y42__R3_BUF_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y43__R0_BUF_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R0_INV_0 (.A(tie_lo_T29Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y43__R1_BUF_0 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R1_INV_0 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R2_INV_0 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y43__R2_INV_1 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y43__R3_BUF_0 (.A(tie_lo_T29Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y44__R0_BUF_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R0_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y44__R1_BUF_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R1_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R2_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y44__R2_INV_1 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y44__R3_BUF_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y45__R0_BUF_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R0_INV_0 (.A(tie_lo_T29Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y45__R1_BUF_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R1_INV_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R2_INV_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y45__R2_INV_1 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y45__R3_BUF_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y46__R0_BUF_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R0_INV_0 (.A(tie_lo_T29Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y46__R1_BUF_0 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R1_INV_0 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R2_INV_0 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y46__R2_INV_1 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y46__R3_BUF_0 (.A(tie_lo_T29Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y47__R0_BUF_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R0_INV_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y47__R1_BUF_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R1_INV_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R2_INV_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y47__R2_INV_1 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y47__R3_BUF_0 (.A(tie_lo_T29Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y48__R0_BUF_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R0_INV_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y48__R1_BUF_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R1_INV_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R2_INV_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y48__R2_INV_1 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y48__R3_BUF_0 (.A(tie_lo_T29Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y49__R0_BUF_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R0_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y49__R1_BUF_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R1_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R2_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y49__R2_INV_1 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y49__R3_BUF_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y4__R0_BUF_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R0_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y4__R1_BUF_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R1_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R2_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y4__R2_INV_1 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y4__R3_BUF_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y50__R0_BUF_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R0_INV_0 (.A(tie_lo_T29Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y50__R1_BUF_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R1_INV_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R2_INV_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y50__R2_INV_1 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y50__R3_BUF_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y51__R0_BUF_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R0_INV_0 (.A(tie_lo_T29Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y51__R1_BUF_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R1_INV_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R2_INV_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y51__R2_INV_1 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y51__R3_BUF_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y52__R0_BUF_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R0_INV_0 (.A(tie_lo_T29Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y52__R1_BUF_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R1_INV_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R2_INV_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y52__R2_INV_1 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y52__R3_BUF_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y53__R0_BUF_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R0_INV_0 (.A(tie_lo_T29Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y53__R1_BUF_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R1_INV_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R2_INV_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y53__R2_INV_1 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y53__R3_BUF_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y54__R0_BUF_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R0_INV_0 (.A(tie_lo_T29Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y54__R1_BUF_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R1_INV_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R2_INV_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y54__R2_INV_1 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y54__R3_BUF_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y55__R0_BUF_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R0_INV_0 (.A(tie_lo_T29Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y55__R1_BUF_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R1_INV_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R2_INV_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y55__R2_INV_1 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y55__R3_BUF_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y56__R0_BUF_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R0_INV_0 (.A(tie_lo_T29Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y56__R1_BUF_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R1_INV_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R2_INV_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y56__R2_INV_1 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y56__R3_BUF_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y57__R0_BUF_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R0_INV_0 (.A(tie_lo_T29Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y57__R1_BUF_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R1_INV_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R2_INV_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y57__R2_INV_1 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y57__R3_BUF_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y58__R0_BUF_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R0_INV_0 (.A(tie_lo_T29Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y58__R1_BUF_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R1_INV_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R2_INV_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y58__R2_INV_1 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y58__R3_BUF_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y59__R0_BUF_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R0_INV_0 (.A(tie_lo_T29Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y59__R1_BUF_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R1_INV_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R2_INV_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y59__R2_INV_1 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y59__R3_BUF_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y5__R0_BUF_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R0_INV_0 (.A(tie_lo_T29Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y5__R1_BUF_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R1_INV_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R2_INV_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y5__R2_INV_1 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y5__R3_BUF_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y60__R0_BUF_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R0_INV_0 (.A(tie_lo_T29Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y60__R1_BUF_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R1_INV_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R2_INV_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y60__R2_INV_1 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y60__R3_BUF_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y61__R0_BUF_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R0_INV_0 (.A(tie_lo_T29Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y61__R1_BUF_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R1_INV_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R2_INV_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y61__R2_INV_1 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y61__R3_BUF_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y62__R0_BUF_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R0_INV_0 (.A(tie_lo_T29Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y62__R1_BUF_0 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R1_INV_0 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R2_INV_0 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y62__R2_INV_1 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y62__R3_BUF_0 (.A(tie_lo_T29Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y63__R0_BUF_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R0_INV_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y63__R1_BUF_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R1_INV_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R2_INV_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y63__R2_INV_1 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y63__R3_BUF_0 (.A(tie_lo_T29Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y64__R0_BUF_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R0_INV_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y64__R1_BUF_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R1_INV_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R2_INV_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y64__R2_INV_1 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y64__R3_BUF_0 (.A(tie_lo_T29Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y65__R0_BUF_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R0_INV_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y65__R1_BUF_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R1_INV_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R2_INV_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y65__R2_INV_1 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y65__R3_BUF_0 (.A(tie_lo_T29Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y66__R0_BUF_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R0_INV_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y66__R1_BUF_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R1_INV_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R2_INV_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y66__R2_INV_1 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y66__R3_BUF_0 (.A(tie_lo_T29Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y67__R0_BUF_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R0_INV_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y67__R1_BUF_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R1_INV_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R2_INV_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y67__R2_INV_1 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y67__R3_BUF_0 (.A(tie_lo_T29Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y68__R0_BUF_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R0_INV_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y68__R1_BUF_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R1_INV_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R2_INV_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y68__R2_INV_1 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y68__R3_BUF_0 (.A(tie_lo_T29Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y69__R0_BUF_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R0_INV_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y69__R1_BUF_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R1_INV_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R2_INV_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y69__R2_INV_1 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y69__R3_BUF_0 (.A(tie_lo_T29Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y6__R0_BUF_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R0_INV_0 (.A(tie_lo_T29Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y6__R1_BUF_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R1_INV_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R2_INV_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y6__R2_INV_1 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y6__R3_BUF_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y70__R0_BUF_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R0_INV_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y70__R1_BUF_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R1_INV_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R2_INV_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y70__R2_INV_1 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y70__R3_BUF_0 (.A(tie_lo_T29Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y71__R0_BUF_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R0_INV_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y71__R1_BUF_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R1_INV_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R2_INV_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y71__R2_INV_1 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y71__R3_BUF_0 (.A(tie_lo_T29Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y72__R0_BUF_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R0_INV_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y72__R1_BUF_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R1_INV_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R2_INV_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y72__R2_INV_1 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y72__R3_BUF_0 (.A(tie_lo_T29Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y73__R0_BUF_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R0_INV_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y73__R1_BUF_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R1_INV_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R2_INV_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y73__R2_INV_1 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y73__R3_BUF_0 (.A(tie_lo_T29Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y74__R0_BUF_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R0_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y74__R1_BUF_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R1_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R2_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y74__R2_INV_1 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y74__R3_BUF_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y75__R0_BUF_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R0_INV_0 (.A(tie_lo_T29Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y75__R1_BUF_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R1_INV_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R2_INV_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y75__R2_INV_1 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y75__R3_BUF_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y76__R0_BUF_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R0_INV_0 (.A(tie_lo_T29Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y76__R1_BUF_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R1_INV_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R2_INV_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y76__R2_INV_1 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y76__R3_BUF_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y77__R0_BUF_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R0_INV_0 (.A(tie_lo_T29Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y77__R1_BUF_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R1_INV_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R2_INV_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y77__R2_INV_1 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y77__R3_BUF_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y78__R0_BUF_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R0_INV_0 (.A(tie_lo_T29Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y78__R1_BUF_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R1_INV_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R2_INV_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y78__R2_INV_1 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y78__R3_BUF_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y79__R0_BUF_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R0_INV_0 (.A(tie_lo_T29Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y79__R1_BUF_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R1_INV_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R2_INV_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y79__R2_INV_1 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y79__R3_BUF_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y7__R0_BUF_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R0_INV_0 (.A(tie_lo_T29Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y7__R1_BUF_0 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R1_INV_0 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R2_INV_0 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y7__R2_INV_1 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y7__R3_BUF_0 (.A(tie_lo_T29Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y80__R0_BUF_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R0_INV_0 (.A(tie_lo_T29Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y80__R1_BUF_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R1_INV_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R2_INV_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y80__R2_INV_1 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y80__R3_BUF_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y81__R0_BUF_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R0_INV_0 (.A(tie_lo_T29Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y81__R1_BUF_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R1_INV_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R2_INV_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y81__R2_INV_1 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y81__R3_BUF_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y82__R0_BUF_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R0_INV_0 (.A(tie_lo_T29Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y82__R1_BUF_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R1_INV_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R2_INV_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y82__R2_INV_1 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y82__R3_BUF_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y83__R0_BUF_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R0_INV_0 (.A(tie_lo_T29Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y83__R1_BUF_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R1_INV_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R2_INV_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y83__R2_INV_1 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y83__R3_BUF_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y84__R0_BUF_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R0_INV_0 (.A(tie_lo_T29Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y84__R1_BUF_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R1_INV_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R2_INV_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y84__R2_INV_1 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y84__R3_BUF_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y85__R0_BUF_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R0_INV_0 (.A(tie_lo_T29Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y85__R1_BUF_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R1_INV_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R2_INV_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y85__R2_INV_1 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y85__R3_BUF_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y86__R0_BUF_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R0_INV_0 (.A(tie_lo_T29Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y86__R1_BUF_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R1_INV_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R2_INV_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y86__R2_INV_1 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y86__R3_BUF_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y87__R0_BUF_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R0_INV_0 (.A(tie_lo_T29Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y87__R1_BUF_0 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R1_INV_0 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R2_INV_0 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y87__R2_INV_1 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y87__R3_BUF_0 (.A(tie_lo_T29Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y88__R0_BUF_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R0_INV_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y88__R1_BUF_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R1_INV_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R2_INV_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y88__R2_INV_1 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y88__R3_BUF_0 (.A(tie_lo_T29Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y89__R0_BUF_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R0_INV_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y89__R1_BUF_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R1_INV_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R2_INV_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y89__R2_INV_1 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y89__R3_BUF_0 (.A(tie_lo_T29Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y8__R0_BUF_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R0_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y8__R1_BUF_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R1_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R2_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y8__R2_INV_1 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y8__R3_BUF_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y9__R0_BUF_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R0_INV_0 (.A(tie_lo_T29Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y9__R1_BUF_0 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R1_INV_0 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T29Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R2_INV_0 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T29Y9__R2_INV_1 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T29Y9__R3_BUF_0 (.A(tie_lo_T29Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y0__R0_BUF_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R0_INV_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y0__R1_BUF_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R1_INV_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R2_INV_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y0__R2_INV_1 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y0__R3_BUF_0 (.A(tie_lo_T2Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y10__R0_BUF_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R0_INV_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y10__R1_BUF_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R1_INV_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R2_INV_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y10__R2_INV_1 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y10__R3_BUF_0 (.A(tie_lo_T2Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y11__R0_BUF_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R0_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y11__R1_BUF_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R1_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R2_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y11__R2_INV_1 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y11__R3_BUF_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y12__R0_BUF_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R0_INV_0 (.A(tie_lo_T2Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y12__R1_BUF_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R1_INV_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R2_INV_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y12__R2_INV_1 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y12__R3_BUF_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y13__R0_BUF_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R0_INV_0 (.A(tie_lo_T2Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y13__R1_BUF_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R1_INV_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R2_INV_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y13__R2_INV_1 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y13__R3_BUF_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y14__R0_BUF_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R0_INV_0 (.A(tie_lo_T2Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y14__R1_BUF_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R1_INV_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R2_INV_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y14__R2_INV_1 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y14__R3_BUF_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y15__R0_BUF_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R0_INV_0 (.A(tie_lo_T2Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y15__R1_BUF_0 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R1_INV_0 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R2_INV_0 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y15__R2_INV_1 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y15__R3_BUF_0 (.A(tie_lo_T2Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y16__R0_BUF_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R0_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y16__R1_BUF_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R1_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R2_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y16__R2_INV_1 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y16__R3_BUF_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y17__R0_BUF_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R0_INV_0 (.A(tie_lo_T2Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y17__R1_BUF_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R1_INV_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R2_INV_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y17__R2_INV_1 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y17__R3_BUF_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y18__R0_BUF_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R0_INV_0 (.A(tie_lo_T2Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y18__R1_BUF_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R1_INV_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R2_INV_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y18__R2_INV_1 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y18__R3_BUF_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y19__R0_BUF_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R0_INV_0 (.A(tie_lo_T2Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y19__R1_BUF_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R1_INV_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R2_INV_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y19__R2_INV_1 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y19__R3_BUF_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y1__R0_BUF_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R0_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y1__R1_BUF_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R1_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R2_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y1__R2_INV_1 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y1__R3_BUF_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y20__R0_BUF_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R0_INV_0 (.A(tie_lo_T2Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y20__R1_BUF_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R1_INV_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R2_INV_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y20__R2_INV_1 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y20__R3_BUF_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y21__R0_BUF_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R0_INV_0 (.A(tie_lo_T2Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y21__R1_BUF_0 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R1_INV_0 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R2_INV_0 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y21__R2_INV_1 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y21__R3_BUF_0 (.A(tie_lo_T2Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y22__R0_BUF_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R0_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y22__R1_BUF_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R1_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R2_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y22__R2_INV_1 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y22__R3_BUF_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y23__R0_BUF_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R0_INV_0 (.A(tie_lo_T2Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y23__R1_BUF_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R1_INV_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R2_INV_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y23__R2_INV_1 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y23__R3_BUF_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y24__R0_BUF_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R0_INV_0 (.A(tie_lo_T2Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y24__R1_BUF_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R1_INV_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R2_INV_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y24__R2_INV_1 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y24__R3_BUF_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y25__R0_BUF_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R0_INV_0 (.A(tie_lo_T2Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y25__R1_BUF_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R1_INV_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R2_INV_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y25__R2_INV_1 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y25__R3_BUF_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y26__R0_BUF_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R0_INV_0 (.A(tie_lo_T2Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y26__R1_BUF_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R1_INV_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R2_INV_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y26__R2_INV_1 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y26__R3_BUF_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y27__R0_BUF_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R0_INV_0 (.A(tie_lo_T2Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y27__R1_BUF_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R1_INV_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R2_INV_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y27__R2_INV_1 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y27__R3_BUF_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y28__R0_BUF_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R0_INV_0 (.A(tie_lo_T2Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y28__R1_BUF_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R1_INV_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R2_INV_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y28__R2_INV_1 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y28__R3_BUF_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y29__R0_BUF_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R0_INV_0 (.A(tie_lo_T2Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y29__R1_BUF_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R1_INV_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R2_INV_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y29__R2_INV_1 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y29__R3_BUF_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y2__R0_BUF_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R0_INV_0 (.A(tie_lo_T2Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y2__R1_BUF_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R1_INV_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R2_INV_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y2__R2_INV_1 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y2__R3_BUF_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y30__R0_BUF_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R0_INV_0 (.A(tie_lo_T2Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y30__R1_BUF_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R1_INV_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R2_INV_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y30__R2_INV_1 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y30__R3_BUF_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y31__R0_BUF_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R0_INV_0 (.A(tie_lo_T2Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y31__R1_BUF_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R1_INV_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R2_INV_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y31__R2_INV_1 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y31__R3_BUF_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y32__R0_BUF_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R0_INV_0 (.A(tie_lo_T2Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y32__R1_BUF_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R1_INV_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R2_INV_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y32__R2_INV_1 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y32__R3_BUF_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y33__R0_BUF_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R0_INV_0 (.A(tie_lo_T2Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y33__R1_BUF_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R1_INV_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R2_INV_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y33__R2_INV_1 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y33__R3_BUF_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y34__R0_BUF_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R0_INV_0 (.A(tie_lo_T2Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y34__R1_BUF_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R1_INV_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R2_INV_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y34__R2_INV_1 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y34__R3_BUF_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y35__R0_BUF_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R0_INV_0 (.A(tie_lo_T2Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y35__R1_BUF_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R1_INV_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R2_INV_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y35__R2_INV_1 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y35__R3_BUF_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y36__R0_BUF_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R0_INV_0 (.A(tie_lo_T2Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y36__R1_BUF_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R1_INV_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R2_INV_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y36__R2_INV_1 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y36__R3_BUF_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y37__R0_BUF_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R0_INV_0 (.A(tie_lo_T2Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y37__R1_BUF_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R1_INV_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R2_INV_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y37__R2_INV_1 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y37__R3_BUF_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y38__R0_BUF_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R0_INV_0 (.A(tie_lo_T2Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y38__R1_BUF_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R1_INV_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R2_INV_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y38__R2_INV_1 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y38__R3_BUF_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y39__R0_BUF_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R0_INV_0 (.A(tie_lo_T2Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y39__R1_BUF_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R1_INV_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R2_INV_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y39__R2_INV_1 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y39__R3_BUF_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y3__R0_BUF_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R0_INV_0 (.A(tie_lo_T2Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y3__R1_BUF_0 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R1_INV_0 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R2_INV_0 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y3__R2_INV_1 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y3__R3_BUF_0 (.A(tie_lo_T2Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y40__R0_BUF_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R0_INV_0 (.A(tie_lo_T2Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y40__R1_BUF_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R1_INV_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R2_INV_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y40__R2_INV_1 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y40__R3_BUF_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y41__R0_BUF_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R0_INV_0 (.A(tie_lo_T2Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y41__R1_BUF_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R1_INV_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R2_INV_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y41__R2_INV_1 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y41__R3_BUF_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y42__R0_BUF_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R0_INV_0 (.A(tie_lo_T2Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y42__R1_BUF_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R1_INV_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R2_INV_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y42__R2_INV_1 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y42__R3_BUF_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y43__R0_BUF_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R0_INV_0 (.A(tie_lo_T2Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y43__R1_BUF_0 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R1_INV_0 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R2_INV_0 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y43__R2_INV_1 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y43__R3_BUF_0 (.A(tie_lo_T2Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y44__R0_BUF_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R0_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y44__R1_BUF_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R1_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R2_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y44__R2_INV_1 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y44__R3_BUF_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y45__R0_BUF_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R0_INV_0 (.A(tie_lo_T2Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y45__R1_BUF_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R1_INV_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R2_INV_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y45__R2_INV_1 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y45__R3_BUF_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y46__R0_BUF_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R0_INV_0 (.A(tie_lo_T2Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y46__R1_BUF_0 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R1_INV_0 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R2_INV_0 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y46__R2_INV_1 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y46__R3_BUF_0 (.A(tie_lo_T2Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y47__R0_BUF_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R0_INV_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y47__R1_BUF_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R1_INV_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R2_INV_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y47__R2_INV_1 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y47__R3_BUF_0 (.A(tie_lo_T2Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y48__R0_BUF_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R0_INV_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y48__R1_BUF_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R1_INV_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R2_INV_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y48__R2_INV_1 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y48__R3_BUF_0 (.A(tie_lo_T2Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y49__R0_BUF_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R0_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y49__R1_BUF_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R1_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R2_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y49__R2_INV_1 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y49__R3_BUF_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y4__R0_BUF_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R0_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y4__R1_BUF_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R1_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R2_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y4__R2_INV_1 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y4__R3_BUF_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y50__R0_BUF_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R0_INV_0 (.A(tie_lo_T2Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y50__R1_BUF_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R1_INV_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R2_INV_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y50__R2_INV_1 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y50__R3_BUF_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y51__R0_BUF_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R0_INV_0 (.A(tie_lo_T2Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y51__R1_BUF_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R1_INV_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R2_INV_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y51__R2_INV_1 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y51__R3_BUF_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y52__R0_BUF_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R0_INV_0 (.A(tie_lo_T2Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y52__R1_BUF_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R1_INV_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R2_INV_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y52__R2_INV_1 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y52__R3_BUF_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y53__R0_BUF_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R0_INV_0 (.A(tie_lo_T2Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y53__R1_BUF_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R1_INV_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R2_INV_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y53__R2_INV_1 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y53__R3_BUF_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y54__R0_BUF_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R0_INV_0 (.A(tie_lo_T2Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y54__R1_BUF_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R1_INV_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R2_INV_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y54__R2_INV_1 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y54__R3_BUF_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y55__R0_BUF_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R0_INV_0 (.A(tie_lo_T2Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y55__R1_BUF_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R1_INV_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R2_INV_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y55__R2_INV_1 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y55__R3_BUF_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y56__R0_BUF_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R0_INV_0 (.A(tie_lo_T2Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y56__R1_BUF_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R1_INV_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R2_INV_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y56__R2_INV_1 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y56__R3_BUF_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y57__R0_BUF_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R0_INV_0 (.A(tie_lo_T2Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y57__R1_BUF_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R1_INV_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R2_INV_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y57__R2_INV_1 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y57__R3_BUF_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y58__R0_BUF_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R0_INV_0 (.A(tie_lo_T2Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y58__R1_BUF_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R1_INV_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R2_INV_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y58__R2_INV_1 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y58__R3_BUF_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y59__R0_BUF_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R0_INV_0 (.A(tie_lo_T2Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y59__R1_BUF_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R1_INV_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R2_INV_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y59__R2_INV_1 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y59__R3_BUF_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y5__R0_BUF_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R0_INV_0 (.A(tie_lo_T2Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y5__R1_BUF_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R1_INV_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R2_INV_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y5__R2_INV_1 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y5__R3_BUF_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y60__R0_BUF_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R0_INV_0 (.A(tie_lo_T2Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y60__R1_BUF_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R1_INV_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R2_INV_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y60__R2_INV_1 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y60__R3_BUF_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y61__R0_BUF_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R0_INV_0 (.A(tie_lo_T2Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y61__R1_BUF_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R1_INV_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R2_INV_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y61__R2_INV_1 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y61__R3_BUF_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y62__R0_BUF_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R0_INV_0 (.A(tie_lo_T2Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y62__R1_BUF_0 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R1_INV_0 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R2_INV_0 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y62__R2_INV_1 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y62__R3_BUF_0 (.A(tie_lo_T2Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y63__R0_BUF_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R0_INV_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y63__R1_BUF_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R1_INV_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R2_INV_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y63__R2_INV_1 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y63__R3_BUF_0 (.A(tie_lo_T2Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y64__R0_BUF_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R0_INV_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y64__R1_BUF_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R1_INV_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R2_INV_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y64__R2_INV_1 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y64__R3_BUF_0 (.A(tie_lo_T2Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y65__R0_BUF_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R0_INV_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y65__R1_BUF_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R1_INV_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R2_INV_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y65__R2_INV_1 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y65__R3_BUF_0 (.A(tie_lo_T2Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y66__R0_BUF_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R0_INV_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y66__R1_BUF_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R1_INV_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R2_INV_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y66__R2_INV_1 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y66__R3_BUF_0 (.A(tie_lo_T2Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y67__R0_BUF_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R0_INV_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y67__R1_BUF_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R1_INV_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R2_INV_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y67__R2_INV_1 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y67__R3_BUF_0 (.A(tie_lo_T2Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y68__R0_BUF_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R0_INV_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y68__R1_BUF_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R1_INV_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R2_INV_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y68__R2_INV_1 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y68__R3_BUF_0 (.A(tie_lo_T2Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y69__R0_BUF_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R0_INV_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y69__R1_BUF_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R1_INV_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R2_INV_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y69__R2_INV_1 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y69__R3_BUF_0 (.A(tie_lo_T2Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y6__R0_BUF_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R0_INV_0 (.A(tie_lo_T2Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y6__R1_BUF_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R1_INV_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R2_INV_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y6__R2_INV_1 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y6__R3_BUF_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y70__R0_BUF_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R0_INV_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y70__R1_BUF_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R1_INV_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R2_INV_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y70__R2_INV_1 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y70__R3_BUF_0 (.A(tie_lo_T2Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y71__R0_BUF_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R0_INV_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y71__R1_BUF_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R1_INV_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R2_INV_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y71__R2_INV_1 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y71__R3_BUF_0 (.A(tie_lo_T2Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y72__R0_BUF_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R0_INV_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y72__R1_BUF_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R1_INV_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R2_INV_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y72__R2_INV_1 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y72__R3_BUF_0 (.A(tie_lo_T2Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y73__R0_BUF_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R0_INV_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y73__R1_BUF_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R1_INV_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R2_INV_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y73__R2_INV_1 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y73__R3_BUF_0 (.A(tie_lo_T2Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y74__R0_BUF_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R0_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y74__R1_BUF_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R1_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R2_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y74__R2_INV_1 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y74__R3_BUF_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y75__R0_BUF_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R0_INV_0 (.A(tie_lo_T2Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y75__R1_BUF_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R1_INV_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R2_INV_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y75__R2_INV_1 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y75__R3_BUF_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y76__R0_BUF_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R0_INV_0 (.A(tie_lo_T2Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y76__R1_BUF_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R1_INV_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R2_INV_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y76__R2_INV_1 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y76__R3_BUF_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y77__R0_BUF_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R0_INV_0 (.A(tie_lo_T2Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y77__R1_BUF_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R1_INV_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R2_INV_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y77__R2_INV_1 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y77__R3_BUF_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y78__R0_BUF_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R0_INV_0 (.A(tie_lo_T2Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y78__R1_BUF_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R1_INV_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R2_INV_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y78__R2_INV_1 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y78__R3_BUF_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y79__R0_BUF_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R0_INV_0 (.A(tie_lo_T2Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y79__R1_BUF_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R1_INV_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R2_INV_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y79__R2_INV_1 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y79__R3_BUF_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y7__R0_BUF_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R0_INV_0 (.A(tie_lo_T2Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y7__R1_BUF_0 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R1_INV_0 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R2_INV_0 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y7__R2_INV_1 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y7__R3_BUF_0 (.A(tie_lo_T2Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y80__R0_BUF_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R0_INV_0 (.A(tie_lo_T2Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y80__R1_BUF_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R1_INV_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R2_INV_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y80__R2_INV_1 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y80__R3_BUF_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y81__R0_BUF_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R0_INV_0 (.A(tie_lo_T2Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y81__R1_BUF_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R1_INV_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R2_INV_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y81__R2_INV_1 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y81__R3_BUF_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y82__R0_BUF_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R0_INV_0 (.A(tie_lo_T2Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y82__R1_BUF_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R1_INV_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R2_INV_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y82__R2_INV_1 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y82__R3_BUF_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y83__R0_BUF_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R0_INV_0 (.A(tie_lo_T2Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y83__R1_BUF_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R1_INV_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R2_INV_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y83__R2_INV_1 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y83__R3_BUF_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y84__R0_BUF_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R0_INV_0 (.A(tie_lo_T2Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y84__R1_BUF_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R1_INV_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R2_INV_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y84__R2_INV_1 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y84__R3_BUF_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y85__R0_BUF_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R0_INV_0 (.A(tie_lo_T2Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y85__R1_BUF_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R1_INV_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R2_INV_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y85__R2_INV_1 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y85__R3_BUF_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y86__R0_BUF_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R0_INV_0 (.A(tie_lo_T2Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y86__R1_BUF_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R1_INV_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R2_INV_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y86__R2_INV_1 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y86__R3_BUF_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y87__R0_BUF_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R0_INV_0 (.A(tie_lo_T2Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y87__R1_BUF_0 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R1_INV_0 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R2_INV_0 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y87__R2_INV_1 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y87__R3_BUF_0 (.A(tie_lo_T2Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y88__R0_BUF_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R0_INV_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y88__R1_BUF_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R1_INV_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R2_INV_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y88__R2_INV_1 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y88__R3_BUF_0 (.A(tie_lo_T2Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y89__R0_BUF_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R0_INV_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y89__R1_BUF_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R1_INV_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R2_INV_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y89__R2_INV_1 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y89__R3_BUF_0 (.A(tie_lo_T2Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y8__R0_BUF_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R0_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y8__R1_BUF_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R1_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R2_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y8__R2_INV_1 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y8__R3_BUF_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y9__R0_BUF_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R0_INV_0 (.A(tie_lo_T2Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y9__R1_BUF_0 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R1_INV_0 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T2Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R2_INV_0 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T2Y9__R2_INV_1 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T2Y9__R3_BUF_0 (.A(tie_lo_T2Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y0__R0_BUF_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R0_INV_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y0__R1_BUF_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R1_INV_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R2_INV_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y0__R2_INV_1 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y0__R3_BUF_0 (.A(tie_lo_T30Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y10__R0_BUF_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R0_INV_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y10__R1_BUF_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R1_INV_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R2_INV_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y10__R2_INV_1 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y10__R3_BUF_0 (.A(tie_lo_T30Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y11__R0_BUF_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R0_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y11__R1_BUF_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R1_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R2_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y11__R2_INV_1 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y11__R3_BUF_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y12__R0_BUF_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R0_INV_0 (.A(tie_lo_T30Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y12__R1_BUF_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R1_INV_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R2_INV_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y12__R2_INV_1 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y12__R3_BUF_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y13__R0_BUF_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R0_INV_0 (.A(tie_lo_T30Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y13__R1_BUF_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R1_INV_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R2_INV_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y13__R2_INV_1 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y13__R3_BUF_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y14__R0_BUF_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R0_INV_0 (.A(tie_lo_T30Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y14__R1_BUF_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R1_INV_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R2_INV_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y14__R2_INV_1 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y14__R3_BUF_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y15__R0_BUF_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R0_INV_0 (.A(tie_lo_T30Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y15__R1_BUF_0 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R1_INV_0 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R2_INV_0 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y15__R2_INV_1 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y15__R3_BUF_0 (.A(tie_lo_T30Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y16__R0_BUF_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R0_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y16__R1_BUF_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R1_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R2_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y16__R2_INV_1 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y16__R3_BUF_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y17__R0_BUF_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R0_INV_0 (.A(tie_lo_T30Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y17__R1_BUF_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R1_INV_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R2_INV_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y17__R2_INV_1 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y17__R3_BUF_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y18__R0_BUF_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R0_INV_0 (.A(tie_lo_T30Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y18__R1_BUF_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R1_INV_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R2_INV_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y18__R2_INV_1 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y18__R3_BUF_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y19__R0_BUF_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R0_INV_0 (.A(tie_lo_T30Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y19__R1_BUF_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R1_INV_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R2_INV_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y19__R2_INV_1 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y19__R3_BUF_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y1__R0_BUF_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R0_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y1__R1_BUF_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R1_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R2_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y1__R2_INV_1 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y1__R3_BUF_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y20__R0_BUF_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R0_INV_0 (.A(tie_lo_T30Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y20__R1_BUF_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R1_INV_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R2_INV_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y20__R2_INV_1 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y20__R3_BUF_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y21__R0_BUF_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R0_INV_0 (.A(tie_lo_T30Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y21__R1_BUF_0 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R1_INV_0 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R2_INV_0 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y21__R2_INV_1 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y21__R3_BUF_0 (.A(tie_lo_T30Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y22__R0_BUF_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R0_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y22__R1_BUF_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R1_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R2_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y22__R2_INV_1 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y22__R3_BUF_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y23__R0_BUF_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R0_INV_0 (.A(tie_lo_T30Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y23__R1_BUF_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R1_INV_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R2_INV_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y23__R2_INV_1 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y23__R3_BUF_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y24__R0_BUF_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R0_INV_0 (.A(tie_lo_T30Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y24__R1_BUF_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R1_INV_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R2_INV_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y24__R2_INV_1 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y24__R3_BUF_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y25__R0_BUF_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R0_INV_0 (.A(tie_lo_T30Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y25__R1_BUF_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R1_INV_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R2_INV_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y25__R2_INV_1 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y25__R3_BUF_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y26__R0_BUF_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R0_INV_0 (.A(tie_lo_T30Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y26__R1_BUF_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R1_INV_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R2_INV_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y26__R2_INV_1 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y26__R3_BUF_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y27__R0_BUF_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R0_INV_0 (.A(tie_lo_T30Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y27__R1_BUF_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R1_INV_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R2_INV_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y27__R2_INV_1 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y27__R3_BUF_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y28__R0_BUF_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R0_INV_0 (.A(tie_lo_T30Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y28__R1_BUF_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R1_INV_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R2_INV_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y28__R2_INV_1 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y28__R3_BUF_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y29__R0_BUF_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R0_INV_0 (.A(tie_lo_T30Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y29__R1_BUF_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R1_INV_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R2_INV_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y29__R2_INV_1 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y29__R3_BUF_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y2__R0_BUF_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R0_INV_0 (.A(tie_lo_T30Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y2__R1_BUF_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R1_INV_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R2_INV_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y2__R2_INV_1 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y2__R3_BUF_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y30__R0_BUF_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R0_INV_0 (.A(tie_lo_T30Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y30__R1_BUF_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R1_INV_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R2_INV_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y30__R2_INV_1 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y30__R3_BUF_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y31__R0_BUF_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R0_INV_0 (.A(tie_lo_T30Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y31__R1_BUF_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R1_INV_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R2_INV_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y31__R2_INV_1 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y31__R3_BUF_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y32__R0_BUF_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R0_INV_0 (.A(tie_lo_T30Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y32__R1_BUF_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R1_INV_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R2_INV_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y32__R2_INV_1 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y32__R3_BUF_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y33__R0_BUF_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R0_INV_0 (.A(tie_lo_T30Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y33__R1_BUF_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R1_INV_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R2_INV_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y33__R2_INV_1 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y33__R3_BUF_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y34__R0_BUF_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R0_INV_0 (.A(tie_lo_T30Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y34__R1_BUF_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R1_INV_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R2_INV_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y34__R2_INV_1 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y34__R3_BUF_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y35__R0_BUF_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R0_INV_0 (.A(tie_lo_T30Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y35__R1_BUF_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R1_INV_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R2_INV_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y35__R2_INV_1 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y35__R3_BUF_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y36__R0_BUF_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R0_INV_0 (.A(tie_lo_T30Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y36__R1_BUF_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R1_INV_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R2_INV_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y36__R2_INV_1 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y36__R3_BUF_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y37__R0_BUF_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R0_INV_0 (.A(tie_lo_T30Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y37__R1_BUF_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R1_INV_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R2_INV_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y37__R2_INV_1 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y37__R3_BUF_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y38__R0_BUF_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R0_INV_0 (.A(tie_lo_T30Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y38__R1_BUF_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R1_INV_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R2_INV_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y38__R2_INV_1 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y38__R3_BUF_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y39__R0_BUF_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R0_INV_0 (.A(tie_lo_T30Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y39__R1_BUF_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R1_INV_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R2_INV_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y39__R2_INV_1 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y39__R3_BUF_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y3__R0_BUF_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R0_INV_0 (.A(tie_lo_T30Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y3__R1_BUF_0 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R1_INV_0 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R2_INV_0 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y3__R2_INV_1 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y3__R3_BUF_0 (.A(tie_lo_T30Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y40__R0_BUF_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R0_INV_0 (.A(tie_lo_T30Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y40__R1_BUF_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R1_INV_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R2_INV_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y40__R2_INV_1 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y40__R3_BUF_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y41__R0_BUF_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R0_INV_0 (.A(tie_lo_T30Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y41__R1_BUF_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R1_INV_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R2_INV_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y41__R2_INV_1 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y41__R3_BUF_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y42__R0_BUF_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R0_INV_0 (.A(tie_lo_T30Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y42__R1_BUF_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R1_INV_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R2_INV_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y42__R2_INV_1 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y42__R3_BUF_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y43__R0_BUF_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R0_INV_0 (.A(tie_lo_T30Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y43__R1_BUF_0 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R1_INV_0 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R2_INV_0 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y43__R2_INV_1 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y43__R3_BUF_0 (.A(tie_lo_T30Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y44__R0_BUF_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R0_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y44__R1_BUF_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R1_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R2_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y44__R2_INV_1 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y44__R3_BUF_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y45__R0_BUF_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R0_INV_0 (.A(tie_lo_T30Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y45__R1_BUF_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R1_INV_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R2_INV_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y45__R2_INV_1 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y45__R3_BUF_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y46__R0_BUF_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R0_INV_0 (.A(tie_lo_T30Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y46__R1_BUF_0 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R1_INV_0 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R2_INV_0 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y46__R2_INV_1 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y46__R3_BUF_0 (.A(tie_lo_T30Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y47__R0_BUF_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R0_INV_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y47__R1_BUF_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R1_INV_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R2_INV_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y47__R2_INV_1 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y47__R3_BUF_0 (.A(tie_lo_T30Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y48__R0_BUF_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R0_INV_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y48__R1_BUF_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R1_INV_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R2_INV_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y48__R2_INV_1 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y48__R3_BUF_0 (.A(tie_lo_T30Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y49__R0_BUF_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R0_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y49__R1_BUF_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R1_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R2_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y49__R2_INV_1 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y49__R3_BUF_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y4__R0_BUF_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R0_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y4__R1_BUF_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R1_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R2_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y4__R2_INV_1 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y4__R3_BUF_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y50__R0_BUF_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R0_INV_0 (.A(tie_lo_T30Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y50__R1_BUF_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R1_INV_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R2_INV_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y50__R2_INV_1 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y50__R3_BUF_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y51__R0_BUF_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R0_INV_0 (.A(tie_lo_T30Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y51__R1_BUF_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R1_INV_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R2_INV_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y51__R2_INV_1 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y51__R3_BUF_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y52__R0_BUF_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R0_INV_0 (.A(tie_lo_T30Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y52__R1_BUF_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R1_INV_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R2_INV_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y52__R2_INV_1 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y52__R3_BUF_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y53__R0_BUF_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R0_INV_0 (.A(tie_lo_T30Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y53__R1_BUF_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R1_INV_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R2_INV_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y53__R2_INV_1 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y53__R3_BUF_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y54__R0_BUF_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R0_INV_0 (.A(tie_lo_T30Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y54__R1_BUF_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R1_INV_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R2_INV_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y54__R2_INV_1 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y54__R3_BUF_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y55__R0_BUF_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R0_INV_0 (.A(tie_lo_T30Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y55__R1_BUF_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R1_INV_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R2_INV_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y55__R2_INV_1 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y55__R3_BUF_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y56__R0_BUF_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R0_INV_0 (.A(tie_lo_T30Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y56__R1_BUF_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R1_INV_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R2_INV_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y56__R2_INV_1 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y56__R3_BUF_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y57__R0_BUF_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R0_INV_0 (.A(tie_lo_T30Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y57__R1_BUF_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R1_INV_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R2_INV_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y57__R2_INV_1 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y57__R3_BUF_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y58__R0_BUF_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R0_INV_0 (.A(tie_lo_T30Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y58__R1_BUF_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R1_INV_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R2_INV_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y58__R2_INV_1 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y58__R3_BUF_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y59__R0_BUF_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R0_INV_0 (.A(tie_lo_T30Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y59__R1_BUF_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R1_INV_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R2_INV_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y59__R2_INV_1 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y59__R3_BUF_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y5__R0_BUF_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R0_INV_0 (.A(tie_lo_T30Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y5__R1_BUF_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R1_INV_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R2_INV_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y5__R2_INV_1 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y5__R3_BUF_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y60__R0_BUF_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R0_INV_0 (.A(tie_lo_T30Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y60__R1_BUF_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R1_INV_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R2_INV_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y60__R2_INV_1 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y60__R3_BUF_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y61__R0_BUF_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R0_INV_0 (.A(tie_lo_T30Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y61__R1_BUF_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R1_INV_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R2_INV_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y61__R2_INV_1 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y61__R3_BUF_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y62__R0_BUF_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R0_INV_0 (.A(tie_lo_T30Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y62__R1_BUF_0 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R1_INV_0 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R2_INV_0 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y62__R2_INV_1 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y62__R3_BUF_0 (.A(tie_lo_T30Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y63__R0_BUF_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R0_INV_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y63__R1_BUF_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R1_INV_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R2_INV_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y63__R2_INV_1 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y63__R3_BUF_0 (.A(tie_lo_T30Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y64__R0_BUF_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R0_INV_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y64__R1_BUF_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R1_INV_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R2_INV_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y64__R2_INV_1 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y64__R3_BUF_0 (.A(tie_lo_T30Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y65__R0_BUF_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R0_INV_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y65__R1_BUF_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R1_INV_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R2_INV_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y65__R2_INV_1 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y65__R3_BUF_0 (.A(tie_lo_T30Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y66__R0_BUF_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R0_INV_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y66__R1_BUF_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R1_INV_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R2_INV_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y66__R2_INV_1 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y66__R3_BUF_0 (.A(tie_lo_T30Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y67__R0_BUF_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R0_INV_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y67__R1_BUF_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R1_INV_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R2_INV_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y67__R2_INV_1 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y67__R3_BUF_0 (.A(tie_lo_T30Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y68__R0_BUF_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R0_INV_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y68__R1_BUF_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R1_INV_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R2_INV_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y68__R2_INV_1 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y68__R3_BUF_0 (.A(tie_lo_T30Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y69__R0_BUF_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R0_INV_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y69__R1_BUF_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R1_INV_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R2_INV_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y69__R2_INV_1 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y69__R3_BUF_0 (.A(tie_lo_T30Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y6__R0_BUF_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R0_INV_0 (.A(tie_lo_T30Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y6__R1_BUF_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R1_INV_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R2_INV_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y6__R2_INV_1 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y6__R3_BUF_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y70__R0_BUF_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R0_INV_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y70__R1_BUF_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R1_INV_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R2_INV_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y70__R2_INV_1 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y70__R3_BUF_0 (.A(tie_lo_T30Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y71__R0_BUF_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R0_INV_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y71__R1_BUF_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R1_INV_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R2_INV_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y71__R2_INV_1 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y71__R3_BUF_0 (.A(tie_lo_T30Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y72__R0_BUF_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R0_INV_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y72__R1_BUF_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R1_INV_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R2_INV_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y72__R2_INV_1 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y72__R3_BUF_0 (.A(tie_lo_T30Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y73__R0_BUF_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R0_INV_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y73__R1_BUF_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R1_INV_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R2_INV_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y73__R2_INV_1 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y73__R3_BUF_0 (.A(tie_lo_T30Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y74__R0_BUF_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R0_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y74__R1_BUF_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R1_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R2_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y74__R2_INV_1 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y74__R3_BUF_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y75__R0_BUF_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R0_INV_0 (.A(tie_lo_T30Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y75__R1_BUF_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R1_INV_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R2_INV_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y75__R2_INV_1 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y75__R3_BUF_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y76__R0_BUF_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R0_INV_0 (.A(tie_lo_T30Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y76__R1_BUF_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R1_INV_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R2_INV_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y76__R2_INV_1 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y76__R3_BUF_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y77__R0_BUF_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R0_INV_0 (.A(tie_lo_T30Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y77__R1_BUF_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R1_INV_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R2_INV_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y77__R2_INV_1 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y77__R3_BUF_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y78__R0_BUF_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R0_INV_0 (.A(tie_lo_T30Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y78__R1_BUF_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R1_INV_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R2_INV_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y78__R2_INV_1 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y78__R3_BUF_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y79__R0_BUF_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R0_INV_0 (.A(tie_lo_T30Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y79__R1_BUF_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R1_INV_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R2_INV_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y79__R2_INV_1 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y79__R3_BUF_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y7__R0_BUF_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R0_INV_0 (.A(tie_lo_T30Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y7__R1_BUF_0 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R1_INV_0 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R2_INV_0 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y7__R2_INV_1 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y7__R3_BUF_0 (.A(tie_lo_T30Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y80__R0_BUF_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R0_INV_0 (.A(tie_lo_T30Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y80__R1_BUF_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R1_INV_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R2_INV_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y80__R2_INV_1 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y80__R3_BUF_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y81__R0_BUF_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R0_INV_0 (.A(tie_lo_T30Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y81__R1_BUF_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R1_INV_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R2_INV_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y81__R2_INV_1 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y81__R3_BUF_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y82__R0_BUF_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R0_INV_0 (.A(tie_lo_T30Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y82__R1_BUF_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R1_INV_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R2_INV_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y82__R2_INV_1 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y82__R3_BUF_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y83__R0_BUF_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R0_INV_0 (.A(tie_lo_T30Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y83__R1_BUF_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R1_INV_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R2_INV_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y83__R2_INV_1 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y83__R3_BUF_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y84__R0_BUF_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R0_INV_0 (.A(tie_lo_T30Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y84__R1_BUF_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R1_INV_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R2_INV_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y84__R2_INV_1 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y84__R3_BUF_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y85__R0_BUF_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R0_INV_0 (.A(tie_lo_T30Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y85__R1_BUF_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R1_INV_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R2_INV_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y85__R2_INV_1 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y85__R3_BUF_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y86__R0_BUF_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R0_INV_0 (.A(tie_lo_T30Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y86__R1_BUF_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R1_INV_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R2_INV_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y86__R2_INV_1 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y86__R3_BUF_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y87__R0_BUF_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R0_INV_0 (.A(tie_lo_T30Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y87__R1_BUF_0 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R1_INV_0 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R2_INV_0 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y87__R2_INV_1 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y87__R3_BUF_0 (.A(tie_lo_T30Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y88__R0_BUF_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R0_INV_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y88__R1_BUF_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R1_INV_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R2_INV_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y88__R2_INV_1 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y88__R3_BUF_0 (.A(tie_lo_T30Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y89__R0_BUF_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R0_INV_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y89__R1_BUF_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R1_INV_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R2_INV_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y89__R2_INV_1 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y89__R3_BUF_0 (.A(tie_lo_T30Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y8__R0_BUF_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R0_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y8__R1_BUF_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R1_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R2_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y8__R2_INV_1 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y8__R3_BUF_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y9__R0_BUF_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R0_INV_0 (.A(tie_lo_T30Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y9__R1_BUF_0 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R1_INV_0 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T30Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R2_INV_0 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T30Y9__R2_INV_1 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T30Y9__R3_BUF_0 (.A(tie_lo_T30Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y0__R0_BUF_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R0_INV_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y0__R1_BUF_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R1_INV_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R2_INV_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y0__R2_INV_1 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y0__R3_BUF_0 (.A(tie_lo_T31Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y10__R0_BUF_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R0_INV_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y10__R1_BUF_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R1_INV_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R2_INV_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y10__R2_INV_1 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y10__R3_BUF_0 (.A(tie_lo_T31Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y11__R0_BUF_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R0_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y11__R1_BUF_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R1_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R2_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y11__R2_INV_1 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y11__R3_BUF_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y12__R0_BUF_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R0_INV_0 (.A(tie_lo_T31Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y12__R1_BUF_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R1_INV_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R2_INV_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y12__R2_INV_1 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y12__R3_BUF_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y13__R0_BUF_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R0_INV_0 (.A(tie_lo_T31Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y13__R1_BUF_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R1_INV_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R2_INV_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y13__R2_INV_1 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y13__R3_BUF_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y14__R0_BUF_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R0_INV_0 (.A(tie_lo_T31Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y14__R1_BUF_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R1_INV_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R2_INV_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y14__R2_INV_1 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y14__R3_BUF_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y15__R0_BUF_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R0_INV_0 (.A(tie_lo_T31Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y15__R1_BUF_0 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R1_INV_0 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R2_INV_0 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y15__R2_INV_1 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y15__R3_BUF_0 (.A(tie_lo_T31Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y16__R0_BUF_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R0_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y16__R1_BUF_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R1_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R2_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y16__R2_INV_1 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y16__R3_BUF_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y17__R0_BUF_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R0_INV_0 (.A(tie_lo_T31Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y17__R1_BUF_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R1_INV_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R2_INV_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y17__R2_INV_1 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y17__R3_BUF_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y18__R0_BUF_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R0_INV_0 (.A(tie_lo_T31Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y18__R1_BUF_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R1_INV_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R2_INV_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y18__R2_INV_1 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y18__R3_BUF_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y19__R0_BUF_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R0_INV_0 (.A(tie_lo_T31Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y19__R1_BUF_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R1_INV_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R2_INV_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y19__R2_INV_1 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y19__R3_BUF_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y1__R0_BUF_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R0_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y1__R1_BUF_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R1_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R2_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y1__R2_INV_1 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y1__R3_BUF_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y20__R0_BUF_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R0_INV_0 (.A(tie_lo_T31Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y20__R1_BUF_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R1_INV_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R2_INV_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y20__R2_INV_1 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y20__R3_BUF_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y21__R0_BUF_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R0_INV_0 (.A(tie_lo_T31Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y21__R1_BUF_0 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R1_INV_0 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R2_INV_0 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y21__R2_INV_1 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y21__R3_BUF_0 (.A(tie_lo_T31Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y22__R0_BUF_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R0_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y22__R1_BUF_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R1_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R2_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y22__R2_INV_1 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y22__R3_BUF_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y23__R0_BUF_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R0_INV_0 (.A(tie_lo_T31Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y23__R1_BUF_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R1_INV_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R2_INV_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y23__R2_INV_1 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y23__R3_BUF_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y24__R0_BUF_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R0_INV_0 (.A(tie_lo_T31Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y24__R1_BUF_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R1_INV_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R2_INV_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y24__R2_INV_1 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y24__R3_BUF_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y25__R0_BUF_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R0_INV_0 (.A(tie_lo_T31Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y25__R1_BUF_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R1_INV_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R2_INV_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y25__R2_INV_1 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y25__R3_BUF_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y26__R0_BUF_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R0_INV_0 (.A(tie_lo_T31Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y26__R1_BUF_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R1_INV_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R2_INV_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y26__R2_INV_1 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y26__R3_BUF_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y27__R0_BUF_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R0_INV_0 (.A(tie_lo_T31Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y27__R1_BUF_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R1_INV_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R2_INV_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y27__R2_INV_1 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y27__R3_BUF_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y28__R0_BUF_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R0_INV_0 (.A(tie_lo_T31Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y28__R1_BUF_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R1_INV_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R2_INV_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y28__R2_INV_1 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y28__R3_BUF_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y29__R0_BUF_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R0_INV_0 (.A(tie_lo_T31Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y29__R1_BUF_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R1_INV_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R2_INV_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y29__R2_INV_1 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y29__R3_BUF_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y2__R0_BUF_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R0_INV_0 (.A(tie_lo_T31Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y2__R1_BUF_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R1_INV_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R2_INV_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y2__R2_INV_1 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y2__R3_BUF_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y30__R0_BUF_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R0_INV_0 (.A(tie_lo_T31Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y30__R1_BUF_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R1_INV_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R2_INV_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y30__R2_INV_1 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y30__R3_BUF_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y31__R0_BUF_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R0_INV_0 (.A(tie_lo_T31Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y31__R1_BUF_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R1_INV_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R2_INV_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y31__R2_INV_1 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y31__R3_BUF_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y32__R0_BUF_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R0_INV_0 (.A(tie_lo_T31Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y32__R1_BUF_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R1_INV_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R2_INV_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y32__R2_INV_1 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y32__R3_BUF_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y33__R0_BUF_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R0_INV_0 (.A(tie_lo_T31Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y33__R1_BUF_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R1_INV_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R2_INV_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y33__R2_INV_1 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y33__R3_BUF_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y34__R0_BUF_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R0_INV_0 (.A(tie_lo_T31Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y34__R1_BUF_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R1_INV_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R2_INV_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y34__R2_INV_1 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y34__R3_BUF_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y35__R0_BUF_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R0_INV_0 (.A(tie_lo_T31Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y35__R1_BUF_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R1_INV_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R2_INV_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y35__R2_INV_1 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y35__R3_BUF_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y36__R0_BUF_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R0_INV_0 (.A(tie_lo_T31Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y36__R1_BUF_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R1_INV_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R2_INV_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y36__R2_INV_1 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y36__R3_BUF_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y37__R0_BUF_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R0_INV_0 (.A(tie_lo_T31Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y37__R1_BUF_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R1_INV_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R2_INV_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y37__R2_INV_1 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y37__R3_BUF_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y38__R0_BUF_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R0_INV_0 (.A(tie_lo_T31Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y38__R1_BUF_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R1_INV_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R2_INV_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y38__R2_INV_1 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y38__R3_BUF_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y39__R0_BUF_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R0_INV_0 (.A(tie_lo_T31Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y39__R1_BUF_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R1_INV_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R2_INV_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y39__R2_INV_1 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y39__R3_BUF_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y3__R0_BUF_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R0_INV_0 (.A(tie_lo_T31Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y3__R1_BUF_0 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R1_INV_0 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R2_INV_0 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y3__R2_INV_1 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y3__R3_BUF_0 (.A(tie_lo_T31Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y40__R0_BUF_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R0_INV_0 (.A(tie_lo_T31Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y40__R1_BUF_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R1_INV_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R2_INV_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y40__R2_INV_1 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y40__R3_BUF_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y41__R0_BUF_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R0_INV_0 (.A(tie_lo_T31Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y41__R1_BUF_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R1_INV_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R2_INV_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y41__R2_INV_1 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y41__R3_BUF_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y42__R0_BUF_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R0_INV_0 (.A(tie_lo_T31Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y42__R1_BUF_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R1_INV_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R2_INV_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y42__R2_INV_1 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y42__R3_BUF_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y43__R0_BUF_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R0_INV_0 (.A(tie_lo_T31Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y43__R1_BUF_0 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R1_INV_0 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R2_INV_0 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y43__R2_INV_1 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y43__R3_BUF_0 (.A(tie_lo_T31Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y44__R0_BUF_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R0_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y44__R1_BUF_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R1_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R2_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y44__R2_INV_1 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y44__R3_BUF_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y45__R0_BUF_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R0_INV_0 (.A(tie_lo_T31Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y45__R1_BUF_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R1_INV_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R2_INV_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y45__R2_INV_1 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y45__R3_BUF_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y46__R0_BUF_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R0_INV_0 (.A(tie_lo_T31Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y46__R1_BUF_0 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R1_INV_0 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R2_INV_0 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y46__R2_INV_1 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y46__R3_BUF_0 (.A(tie_lo_T31Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y47__R0_BUF_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R0_INV_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y47__R1_BUF_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R1_INV_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R2_INV_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y47__R2_INV_1 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y47__R3_BUF_0 (.A(tie_lo_T31Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y48__R0_BUF_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R0_INV_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y48__R1_BUF_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R1_INV_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R2_INV_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y48__R2_INV_1 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y48__R3_BUF_0 (.A(tie_lo_T31Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y49__R0_BUF_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R0_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y49__R1_BUF_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R1_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R2_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y49__R2_INV_1 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y49__R3_BUF_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y4__R0_BUF_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R0_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y4__R1_BUF_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R1_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R2_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y4__R2_INV_1 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y4__R3_BUF_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y50__R0_BUF_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R0_INV_0 (.A(tie_lo_T31Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y50__R1_BUF_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R1_INV_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R2_INV_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y50__R2_INV_1 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y50__R3_BUF_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y51__R0_BUF_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R0_INV_0 (.A(tie_lo_T31Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y51__R1_BUF_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R1_INV_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R2_INV_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y51__R2_INV_1 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y51__R3_BUF_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y52__R0_BUF_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R0_INV_0 (.A(tie_lo_T31Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y52__R1_BUF_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R1_INV_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R2_INV_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y52__R2_INV_1 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y52__R3_BUF_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y53__R0_BUF_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R0_INV_0 (.A(tie_lo_T31Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y53__R1_BUF_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R1_INV_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R2_INV_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y53__R2_INV_1 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y53__R3_BUF_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y54__R0_BUF_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R0_INV_0 (.A(tie_lo_T31Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y54__R1_BUF_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R1_INV_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R2_INV_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y54__R2_INV_1 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y54__R3_BUF_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y55__R0_BUF_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R0_INV_0 (.A(tie_lo_T31Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y55__R1_BUF_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R1_INV_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R2_INV_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y55__R2_INV_1 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y55__R3_BUF_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y56__R0_BUF_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R0_INV_0 (.A(tie_lo_T31Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y56__R1_BUF_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R1_INV_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R2_INV_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y56__R2_INV_1 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y56__R3_BUF_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y57__R0_BUF_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R0_INV_0 (.A(tie_lo_T31Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y57__R1_BUF_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R1_INV_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R2_INV_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y57__R2_INV_1 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y57__R3_BUF_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y58__R0_BUF_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R0_INV_0 (.A(tie_lo_T31Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y58__R1_BUF_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R1_INV_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R2_INV_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y58__R2_INV_1 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y58__R3_BUF_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y59__R0_BUF_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R0_INV_0 (.A(tie_lo_T31Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y59__R1_BUF_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R1_INV_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R2_INV_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y59__R2_INV_1 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y59__R3_BUF_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y5__R0_BUF_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R0_INV_0 (.A(tie_lo_T31Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y5__R1_BUF_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R1_INV_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R2_INV_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y5__R2_INV_1 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y5__R3_BUF_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y60__R0_BUF_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R0_INV_0 (.A(tie_lo_T31Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y60__R1_BUF_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R1_INV_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R2_INV_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y60__R2_INV_1 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y60__R3_BUF_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y61__R0_BUF_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R0_INV_0 (.A(tie_lo_T31Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y61__R1_BUF_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R1_INV_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R2_INV_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y61__R2_INV_1 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y61__R3_BUF_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y62__R0_BUF_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R0_INV_0 (.A(tie_lo_T31Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y62__R1_BUF_0 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R1_INV_0 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R2_INV_0 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y62__R2_INV_1 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y62__R3_BUF_0 (.A(tie_lo_T31Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y63__R0_BUF_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R0_INV_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y63__R1_BUF_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R1_INV_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R2_INV_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y63__R2_INV_1 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y63__R3_BUF_0 (.A(tie_lo_T31Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y64__R0_BUF_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R0_INV_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y64__R1_BUF_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R1_INV_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R2_INV_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y64__R2_INV_1 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y64__R3_BUF_0 (.A(tie_lo_T31Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y65__R0_BUF_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R0_INV_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y65__R1_BUF_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R1_INV_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R2_INV_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y65__R2_INV_1 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y65__R3_BUF_0 (.A(tie_lo_T31Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y66__R0_BUF_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R0_INV_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y66__R1_BUF_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R1_INV_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R2_INV_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y66__R2_INV_1 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y66__R3_BUF_0 (.A(tie_lo_T31Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y67__R0_BUF_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R0_INV_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y67__R1_BUF_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R1_INV_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R2_INV_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y67__R2_INV_1 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y67__R3_BUF_0 (.A(tie_lo_T31Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y68__R0_BUF_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R0_INV_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y68__R1_BUF_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R1_INV_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R2_INV_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y68__R2_INV_1 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y68__R3_BUF_0 (.A(tie_lo_T31Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y69__R0_BUF_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R0_INV_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y69__R1_BUF_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R1_INV_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R2_INV_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y69__R2_INV_1 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y69__R3_BUF_0 (.A(tie_lo_T31Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y6__R0_BUF_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R0_INV_0 (.A(tie_lo_T31Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y6__R1_BUF_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R1_INV_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R2_INV_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y6__R2_INV_1 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y6__R3_BUF_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y70__R0_BUF_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R0_INV_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y70__R1_BUF_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R1_INV_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R2_INV_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y70__R2_INV_1 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y70__R3_BUF_0 (.A(tie_lo_T31Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y71__R0_BUF_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R0_INV_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y71__R1_BUF_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R1_INV_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R2_INV_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y71__R2_INV_1 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y71__R3_BUF_0 (.A(tie_lo_T31Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y72__R0_BUF_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R0_INV_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y72__R1_BUF_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R1_INV_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R2_INV_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y72__R2_INV_1 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y72__R3_BUF_0 (.A(tie_lo_T31Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y73__R0_BUF_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R0_INV_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y73__R1_BUF_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R1_INV_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R2_INV_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y73__R2_INV_1 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y73__R3_BUF_0 (.A(tie_lo_T31Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y74__R0_BUF_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R0_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y74__R1_BUF_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R1_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R2_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y74__R2_INV_1 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y74__R3_BUF_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y75__R0_BUF_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R0_INV_0 (.A(tie_lo_T31Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y75__R1_BUF_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R1_INV_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R2_INV_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y75__R2_INV_1 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y75__R3_BUF_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y76__R0_BUF_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R0_INV_0 (.A(tie_lo_T31Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y76__R1_BUF_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R1_INV_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R2_INV_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y76__R2_INV_1 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y76__R3_BUF_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y77__R0_BUF_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R0_INV_0 (.A(tie_lo_T31Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y77__R1_BUF_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R1_INV_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R2_INV_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y77__R2_INV_1 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y77__R3_BUF_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y78__R0_BUF_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R0_INV_0 (.A(tie_lo_T31Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y78__R1_BUF_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R1_INV_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R2_INV_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y78__R2_INV_1 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y78__R3_BUF_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y79__R0_BUF_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R0_INV_0 (.A(tie_lo_T31Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y79__R1_BUF_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R1_INV_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R2_INV_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y79__R2_INV_1 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y79__R3_BUF_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y7__R0_BUF_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R0_INV_0 (.A(tie_lo_T31Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y7__R1_BUF_0 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R1_INV_0 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R2_INV_0 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y7__R2_INV_1 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y7__R3_BUF_0 (.A(tie_lo_T31Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y80__R0_BUF_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R0_INV_0 (.A(tie_lo_T31Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y80__R1_BUF_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R1_INV_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R2_INV_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y80__R2_INV_1 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y80__R3_BUF_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y81__R0_BUF_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R0_INV_0 (.A(tie_lo_T31Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y81__R1_BUF_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R1_INV_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R2_INV_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y81__R2_INV_1 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y81__R3_BUF_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y82__R0_BUF_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R0_INV_0 (.A(tie_lo_T31Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y82__R1_BUF_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R1_INV_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R2_INV_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y82__R2_INV_1 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y82__R3_BUF_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y83__R0_BUF_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R0_INV_0 (.A(tie_lo_T31Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y83__R1_BUF_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R1_INV_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R2_INV_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y83__R2_INV_1 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y83__R3_BUF_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y84__R0_BUF_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R0_INV_0 (.A(tie_lo_T31Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y84__R1_BUF_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R1_INV_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R2_INV_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y84__R2_INV_1 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y84__R3_BUF_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y85__R0_BUF_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R0_INV_0 (.A(tie_lo_T31Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y85__R1_BUF_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R1_INV_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R2_INV_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y85__R2_INV_1 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y85__R3_BUF_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y86__R0_BUF_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R0_INV_0 (.A(tie_lo_T31Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y86__R1_BUF_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R1_INV_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R2_INV_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y86__R2_INV_1 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y86__R3_BUF_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y87__R0_BUF_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R0_INV_0 (.A(tie_lo_T31Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y87__R1_BUF_0 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R1_INV_0 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R2_INV_0 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y87__R2_INV_1 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y87__R3_BUF_0 (.A(tie_lo_T31Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y88__R0_BUF_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R0_INV_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y88__R1_BUF_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R1_INV_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R2_INV_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y88__R2_INV_1 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y88__R3_BUF_0 (.A(tie_lo_T31Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y89__R0_BUF_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R0_INV_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y89__R1_BUF_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R1_INV_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R2_INV_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y89__R2_INV_1 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y89__R3_BUF_0 (.A(tie_lo_T31Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y8__R0_BUF_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R0_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y8__R1_BUF_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R1_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R2_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y8__R2_INV_1 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y8__R3_BUF_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y9__R0_BUF_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R0_INV_0 (.A(tie_lo_T31Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y9__R1_BUF_0 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R1_INV_0 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T31Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R2_INV_0 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T31Y9__R2_INV_1 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T31Y9__R3_BUF_0 (.A(tie_lo_T31Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y0__R0_BUF_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R0_INV_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y0__R1_BUF_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R1_INV_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R2_INV_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y0__R2_INV_1 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y0__R3_BUF_0 (.A(tie_lo_T32Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y10__R0_BUF_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R0_INV_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y10__R1_BUF_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R1_INV_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R2_INV_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y10__R2_INV_1 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y10__R3_BUF_0 (.A(tie_lo_T32Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y11__R0_BUF_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R0_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y11__R1_BUF_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R1_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R2_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y11__R2_INV_1 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y11__R3_BUF_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y12__R0_BUF_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R0_INV_0 (.A(tie_lo_T32Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y12__R1_BUF_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R1_INV_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R2_INV_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y12__R2_INV_1 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y12__R3_BUF_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y13__R0_BUF_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R0_INV_0 (.A(tie_lo_T32Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y13__R1_BUF_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R1_INV_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R2_INV_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y13__R2_INV_1 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y13__R3_BUF_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y14__R0_BUF_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R0_INV_0 (.A(tie_lo_T32Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y14__R1_BUF_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R1_INV_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R2_INV_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y14__R2_INV_1 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y14__R3_BUF_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y15__R0_BUF_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R0_INV_0 (.A(tie_lo_T32Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y15__R1_BUF_0 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R1_INV_0 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R2_INV_0 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y15__R2_INV_1 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y15__R3_BUF_0 (.A(tie_lo_T32Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y16__R0_BUF_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R0_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y16__R1_BUF_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R1_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R2_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y16__R2_INV_1 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y16__R3_BUF_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y17__R0_BUF_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R0_INV_0 (.A(tie_lo_T32Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y17__R1_BUF_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R1_INV_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R2_INV_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y17__R2_INV_1 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y17__R3_BUF_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y18__R0_BUF_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R0_INV_0 (.A(tie_lo_T32Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y18__R1_BUF_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R1_INV_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R2_INV_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y18__R2_INV_1 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y18__R3_BUF_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y19__R0_BUF_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R0_INV_0 (.A(tie_lo_T32Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y19__R1_BUF_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R1_INV_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R2_INV_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y19__R2_INV_1 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y19__R3_BUF_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y1__R0_BUF_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R0_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y1__R1_BUF_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R1_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R2_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y1__R2_INV_1 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y1__R3_BUF_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y20__R0_BUF_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R0_INV_0 (.A(tie_lo_T32Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y20__R1_BUF_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R1_INV_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R2_INV_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y20__R2_INV_1 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y20__R3_BUF_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y21__R0_BUF_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R0_INV_0 (.A(tie_lo_T32Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y21__R1_BUF_0 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R1_INV_0 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R2_INV_0 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y21__R2_INV_1 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y21__R3_BUF_0 (.A(tie_lo_T32Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y22__R0_BUF_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R0_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y22__R1_BUF_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R1_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R2_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y22__R2_INV_1 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y22__R3_BUF_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y23__R0_BUF_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R0_INV_0 (.A(tie_lo_T32Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y23__R1_BUF_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R1_INV_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R2_INV_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y23__R2_INV_1 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y23__R3_BUF_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y24__R0_BUF_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R0_INV_0 (.A(tie_lo_T32Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y24__R1_BUF_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R1_INV_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R2_INV_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y24__R2_INV_1 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y24__R3_BUF_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y25__R0_BUF_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R0_INV_0 (.A(tie_lo_T32Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y25__R1_BUF_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R1_INV_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R2_INV_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y25__R2_INV_1 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y25__R3_BUF_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y26__R0_BUF_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R0_INV_0 (.A(tie_lo_T32Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y26__R1_BUF_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R1_INV_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R2_INV_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y26__R2_INV_1 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y26__R3_BUF_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y27__R0_BUF_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R0_INV_0 (.A(tie_lo_T32Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y27__R1_BUF_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R1_INV_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R2_INV_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y27__R2_INV_1 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y27__R3_BUF_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y28__R0_BUF_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R0_INV_0 (.A(tie_lo_T32Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y28__R1_BUF_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R1_INV_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R2_INV_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y28__R2_INV_1 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y28__R3_BUF_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y29__R0_BUF_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R0_INV_0 (.A(tie_lo_T32Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y29__R1_BUF_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R1_INV_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R2_INV_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y29__R2_INV_1 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y29__R3_BUF_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y2__R0_BUF_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R0_INV_0 (.A(tie_lo_T32Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y2__R1_BUF_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R1_INV_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R2_INV_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y2__R2_INV_1 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y2__R3_BUF_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y30__R0_BUF_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R0_INV_0 (.A(tie_lo_T32Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y30__R1_BUF_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R1_INV_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R2_INV_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y30__R2_INV_1 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y30__R3_BUF_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y31__R0_BUF_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R0_INV_0 (.A(tie_lo_T32Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y31__R1_BUF_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R1_INV_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R2_INV_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y31__R2_INV_1 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y31__R3_BUF_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y32__R0_BUF_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R0_INV_0 (.A(tie_lo_T32Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y32__R1_BUF_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R1_INV_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R2_INV_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y32__R2_INV_1 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y32__R3_BUF_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y33__R0_BUF_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R0_INV_0 (.A(tie_lo_T32Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y33__R1_BUF_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R1_INV_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R2_INV_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y33__R2_INV_1 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y33__R3_BUF_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y34__R0_BUF_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R0_INV_0 (.A(tie_lo_T32Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y34__R1_BUF_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R1_INV_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R2_INV_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y34__R2_INV_1 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y34__R3_BUF_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y35__R0_BUF_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R0_INV_0 (.A(tie_lo_T32Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y35__R1_BUF_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R1_INV_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R2_INV_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y35__R2_INV_1 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y35__R3_BUF_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y36__R0_BUF_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R0_INV_0 (.A(tie_lo_T32Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y36__R1_BUF_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R1_INV_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R2_INV_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y36__R2_INV_1 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y36__R3_BUF_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y37__R0_BUF_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R0_INV_0 (.A(tie_lo_T32Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y37__R1_BUF_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R1_INV_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R2_INV_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y37__R2_INV_1 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y37__R3_BUF_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y38__R0_BUF_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R0_INV_0 (.A(tie_lo_T32Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y38__R1_BUF_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R1_INV_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R2_INV_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y38__R2_INV_1 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y38__R3_BUF_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y39__R0_BUF_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R0_INV_0 (.A(tie_lo_T32Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y39__R1_BUF_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R1_INV_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R2_INV_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y39__R2_INV_1 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y39__R3_BUF_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y3__R0_BUF_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R0_INV_0 (.A(tie_lo_T32Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y3__R1_BUF_0 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R1_INV_0 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R2_INV_0 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y3__R2_INV_1 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y3__R3_BUF_0 (.A(tie_lo_T32Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y40__R0_BUF_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R0_INV_0 (.A(tie_lo_T32Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y40__R1_BUF_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R1_INV_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R2_INV_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y40__R2_INV_1 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y40__R3_BUF_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y41__R0_BUF_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R0_INV_0 (.A(tie_lo_T32Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y41__R1_BUF_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R1_INV_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R2_INV_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y41__R2_INV_1 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y41__R3_BUF_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y42__R0_BUF_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R0_INV_0 (.A(tie_lo_T32Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y42__R1_BUF_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R1_INV_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R2_INV_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y42__R2_INV_1 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y42__R3_BUF_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y43__R0_BUF_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R0_INV_0 (.A(tie_lo_T32Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y43__R1_BUF_0 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R1_INV_0 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R2_INV_0 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y43__R2_INV_1 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y43__R3_BUF_0 (.A(tie_lo_T32Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y44__R0_BUF_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R0_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y44__R1_BUF_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R1_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R2_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y44__R2_INV_1 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y44__R3_BUF_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y45__R0_BUF_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R0_INV_0 (.A(tie_lo_T32Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y45__R1_BUF_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R1_INV_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R2_INV_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y45__R2_INV_1 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y45__R3_BUF_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y46__R0_BUF_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R0_INV_0 (.A(tie_lo_T32Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y46__R1_BUF_0 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R1_INV_0 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R2_INV_0 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y46__R2_INV_1 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y46__R3_BUF_0 (.A(tie_lo_T32Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y47__R0_BUF_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R0_INV_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y47__R1_BUF_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R1_INV_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R2_INV_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y47__R2_INV_1 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y47__R3_BUF_0 (.A(tie_lo_T32Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y48__R0_BUF_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R0_INV_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y48__R1_BUF_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R1_INV_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R2_INV_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y48__R2_INV_1 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y48__R3_BUF_0 (.A(tie_lo_T32Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y49__R0_BUF_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R0_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y49__R1_BUF_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R1_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R2_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y49__R2_INV_1 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y49__R3_BUF_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y4__R0_BUF_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R0_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y4__R1_BUF_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R1_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R2_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y4__R2_INV_1 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y4__R3_BUF_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y50__R0_BUF_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R0_INV_0 (.A(tie_lo_T32Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y50__R1_BUF_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R1_INV_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R2_INV_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y50__R2_INV_1 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y50__R3_BUF_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y51__R0_BUF_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R0_INV_0 (.A(tie_lo_T32Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y51__R1_BUF_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R1_INV_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R2_INV_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y51__R2_INV_1 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y51__R3_BUF_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y52__R0_BUF_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R0_INV_0 (.A(tie_lo_T32Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y52__R1_BUF_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R1_INV_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R2_INV_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y52__R2_INV_1 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y52__R3_BUF_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y53__R0_BUF_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R0_INV_0 (.A(tie_lo_T32Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y53__R1_BUF_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R1_INV_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R2_INV_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y53__R2_INV_1 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y53__R3_BUF_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y54__R0_BUF_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R0_INV_0 (.A(tie_lo_T32Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y54__R1_BUF_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R1_INV_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R2_INV_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y54__R2_INV_1 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y54__R3_BUF_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y55__R0_BUF_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R0_INV_0 (.A(tie_lo_T32Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y55__R1_BUF_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R1_INV_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R2_INV_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y55__R2_INV_1 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y55__R3_BUF_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y56__R0_BUF_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R0_INV_0 (.A(tie_lo_T32Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y56__R1_BUF_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R1_INV_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R2_INV_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y56__R2_INV_1 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y56__R3_BUF_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y57__R0_BUF_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R0_INV_0 (.A(tie_lo_T32Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y57__R1_BUF_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R1_INV_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R2_INV_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y57__R2_INV_1 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y57__R3_BUF_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y58__R0_BUF_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R0_INV_0 (.A(tie_lo_T32Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y58__R1_BUF_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R1_INV_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R2_INV_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y58__R2_INV_1 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y58__R3_BUF_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y59__R0_BUF_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R0_INV_0 (.A(tie_lo_T32Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y59__R1_BUF_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R1_INV_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R2_INV_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y59__R2_INV_1 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y59__R3_BUF_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y5__R0_BUF_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R0_INV_0 (.A(tie_lo_T32Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y5__R1_BUF_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R1_INV_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R2_INV_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y5__R2_INV_1 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y5__R3_BUF_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y60__R0_BUF_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R0_INV_0 (.A(tie_lo_T32Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y60__R1_BUF_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R1_INV_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R2_INV_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y60__R2_INV_1 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y60__R3_BUF_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y61__R0_BUF_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R0_INV_0 (.A(tie_lo_T32Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y61__R1_BUF_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R1_INV_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R2_INV_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y61__R2_INV_1 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y61__R3_BUF_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y62__R0_BUF_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R0_INV_0 (.A(tie_lo_T32Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y62__R1_BUF_0 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R1_INV_0 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R2_INV_0 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y62__R2_INV_1 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y62__R3_BUF_0 (.A(tie_lo_T32Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y63__R0_BUF_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R0_INV_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y63__R1_BUF_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R1_INV_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R2_INV_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y63__R2_INV_1 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y63__R3_BUF_0 (.A(tie_lo_T32Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y64__R0_BUF_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R0_INV_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y64__R1_BUF_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R1_INV_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R2_INV_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y64__R2_INV_1 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y64__R3_BUF_0 (.A(tie_lo_T32Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y65__R0_BUF_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R0_INV_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y65__R1_BUF_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R1_INV_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R2_INV_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y65__R2_INV_1 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y65__R3_BUF_0 (.A(tie_lo_T32Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y66__R0_BUF_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R0_INV_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y66__R1_BUF_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R1_INV_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R2_INV_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y66__R2_INV_1 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y66__R3_BUF_0 (.A(tie_lo_T32Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y67__R0_BUF_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R0_INV_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y67__R1_BUF_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R1_INV_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R2_INV_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y67__R2_INV_1 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y67__R3_BUF_0 (.A(tie_lo_T32Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y68__R0_BUF_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R0_INV_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y68__R1_BUF_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R1_INV_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R2_INV_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y68__R2_INV_1 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y68__R3_BUF_0 (.A(tie_lo_T32Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y69__R0_BUF_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R0_INV_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y69__R1_BUF_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R1_INV_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R2_INV_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y69__R2_INV_1 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y69__R3_BUF_0 (.A(tie_lo_T32Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y6__R0_BUF_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R0_INV_0 (.A(tie_lo_T32Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y6__R1_BUF_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R1_INV_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R2_INV_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y6__R2_INV_1 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y6__R3_BUF_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y70__R0_BUF_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R0_INV_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y70__R1_BUF_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R1_INV_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R2_INV_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y70__R2_INV_1 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y70__R3_BUF_0 (.A(tie_lo_T32Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y71__R0_BUF_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R0_INV_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y71__R1_BUF_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R1_INV_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R2_INV_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y71__R2_INV_1 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y71__R3_BUF_0 (.A(tie_lo_T32Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y72__R0_BUF_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R0_INV_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y72__R1_BUF_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R1_INV_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R2_INV_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y72__R2_INV_1 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y72__R3_BUF_0 (.A(tie_lo_T32Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y73__R0_BUF_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R0_INV_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y73__R1_BUF_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R1_INV_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R2_INV_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y73__R2_INV_1 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y73__R3_BUF_0 (.A(tie_lo_T32Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y74__R0_BUF_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R0_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y74__R1_BUF_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R1_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R2_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y74__R2_INV_1 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y74__R3_BUF_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y75__R0_BUF_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R0_INV_0 (.A(tie_lo_T32Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y75__R1_BUF_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R1_INV_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R2_INV_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y75__R2_INV_1 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y75__R3_BUF_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y76__R0_BUF_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R0_INV_0 (.A(tie_lo_T32Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y76__R1_BUF_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R1_INV_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R2_INV_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y76__R2_INV_1 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y76__R3_BUF_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y77__R0_BUF_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R0_INV_0 (.A(tie_lo_T32Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y77__R1_BUF_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R1_INV_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R2_INV_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y77__R2_INV_1 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y77__R3_BUF_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y78__R0_BUF_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R0_INV_0 (.A(tie_lo_T32Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y78__R1_BUF_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R1_INV_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R2_INV_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y78__R2_INV_1 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y78__R3_BUF_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y79__R0_BUF_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R0_INV_0 (.A(tie_lo_T32Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y79__R1_BUF_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R1_INV_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R2_INV_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y79__R2_INV_1 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y79__R3_BUF_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y7__R0_BUF_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R0_INV_0 (.A(tie_lo_T32Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y7__R1_BUF_0 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R1_INV_0 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R2_INV_0 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y7__R2_INV_1 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y7__R3_BUF_0 (.A(tie_lo_T32Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y80__R0_BUF_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R0_INV_0 (.A(tie_lo_T32Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y80__R1_BUF_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R1_INV_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R2_INV_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y80__R2_INV_1 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y80__R3_BUF_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y81__R0_BUF_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R0_INV_0 (.A(tie_lo_T32Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y81__R1_BUF_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R1_INV_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R2_INV_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y81__R2_INV_1 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y81__R3_BUF_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y82__R0_BUF_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R0_INV_0 (.A(tie_lo_T32Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y82__R1_BUF_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R1_INV_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R2_INV_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y82__R2_INV_1 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y82__R3_BUF_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y83__R0_BUF_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R0_INV_0 (.A(tie_lo_T32Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y83__R1_BUF_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R1_INV_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R2_INV_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y83__R2_INV_1 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y83__R3_BUF_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y84__R0_BUF_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R0_INV_0 (.A(tie_lo_T32Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y84__R1_BUF_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R1_INV_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R2_INV_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y84__R2_INV_1 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y84__R3_BUF_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y85__R0_BUF_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R0_INV_0 (.A(tie_lo_T32Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y85__R1_BUF_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R1_INV_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R2_INV_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y85__R2_INV_1 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y85__R3_BUF_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y86__R0_BUF_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R0_INV_0 (.A(tie_lo_T32Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y86__R1_BUF_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R1_INV_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R2_INV_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y86__R2_INV_1 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y86__R3_BUF_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y87__R0_BUF_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R0_INV_0 (.A(tie_lo_T32Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y87__R1_BUF_0 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R1_INV_0 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R2_INV_0 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y87__R2_INV_1 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y87__R3_BUF_0 (.A(tie_lo_T32Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y88__R0_BUF_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R0_INV_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y88__R1_BUF_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R1_INV_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R2_INV_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y88__R2_INV_1 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y88__R3_BUF_0 (.A(tie_lo_T32Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y89__R0_BUF_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R0_INV_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y89__R1_BUF_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R1_INV_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R2_INV_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y89__R2_INV_1 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y89__R3_BUF_0 (.A(tie_lo_T32Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y8__R0_BUF_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R0_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y8__R1_BUF_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R1_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R2_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y8__R2_INV_1 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y8__R3_BUF_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y9__R0_BUF_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R0_INV_0 (.A(tie_lo_T32Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y9__R1_BUF_0 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R1_INV_0 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T32Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R2_INV_0 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T32Y9__R2_INV_1 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T32Y9__R3_BUF_0 (.A(tie_lo_T32Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y0__R0_BUF_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R0_INV_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y0__R1_BUF_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R1_INV_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R2_INV_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y0__R2_INV_1 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y0__R3_BUF_0 (.A(tie_lo_T33Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y10__R0_BUF_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R0_INV_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y10__R1_BUF_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R1_INV_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R2_INV_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y10__R2_INV_1 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y10__R3_BUF_0 (.A(tie_lo_T33Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y11__R0_BUF_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R0_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y11__R1_BUF_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R1_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R2_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y11__R2_INV_1 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y11__R3_BUF_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y12__R0_BUF_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R0_INV_0 (.A(tie_lo_T33Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y12__R1_BUF_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R1_INV_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R2_INV_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y12__R2_INV_1 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y12__R3_BUF_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y13__R0_BUF_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R0_INV_0 (.A(tie_lo_T33Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y13__R1_BUF_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R1_INV_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R2_INV_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y13__R2_INV_1 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y13__R3_BUF_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y14__R0_BUF_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R0_INV_0 (.A(tie_lo_T33Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y14__R1_BUF_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R1_INV_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R2_INV_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y14__R2_INV_1 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y14__R3_BUF_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y15__R0_BUF_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R0_INV_0 (.A(tie_lo_T33Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y15__R1_BUF_0 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R1_INV_0 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R2_INV_0 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y15__R2_INV_1 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y15__R3_BUF_0 (.A(tie_lo_T33Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y16__R0_BUF_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R0_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y16__R1_BUF_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R1_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R2_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y16__R2_INV_1 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y16__R3_BUF_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y17__R0_BUF_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R0_INV_0 (.A(tie_lo_T33Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y17__R1_BUF_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R1_INV_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R2_INV_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y17__R2_INV_1 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y17__R3_BUF_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y18__R0_BUF_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R0_INV_0 (.A(tie_lo_T33Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y18__R1_BUF_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R1_INV_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R2_INV_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y18__R2_INV_1 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y18__R3_BUF_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y19__R0_BUF_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R0_INV_0 (.A(tie_lo_T33Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y19__R1_BUF_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R1_INV_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R2_INV_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y19__R2_INV_1 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y19__R3_BUF_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y1__R0_BUF_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R0_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y1__R1_BUF_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R1_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R2_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y1__R2_INV_1 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y1__R3_BUF_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y20__R0_BUF_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R0_INV_0 (.A(tie_lo_T33Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y20__R1_BUF_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R1_INV_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R2_INV_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y20__R2_INV_1 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y20__R3_BUF_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y21__R0_BUF_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R0_INV_0 (.A(tie_lo_T33Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y21__R1_BUF_0 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R1_INV_0 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R2_INV_0 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y21__R2_INV_1 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y21__R3_BUF_0 (.A(tie_lo_T33Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y22__R0_BUF_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R0_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y22__R1_BUF_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R1_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R2_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y22__R2_INV_1 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y22__R3_BUF_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y23__R0_BUF_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R0_INV_0 (.A(tie_lo_T33Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y23__R1_BUF_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R1_INV_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R2_INV_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y23__R2_INV_1 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y23__R3_BUF_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y24__R0_BUF_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R0_INV_0 (.A(tie_lo_T33Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y24__R1_BUF_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R1_INV_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R2_INV_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y24__R2_INV_1 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y24__R3_BUF_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y25__R0_BUF_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R0_INV_0 (.A(tie_lo_T33Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y25__R1_BUF_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R1_INV_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R2_INV_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y25__R2_INV_1 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y25__R3_BUF_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y26__R0_BUF_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R0_INV_0 (.A(tie_lo_T33Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y26__R1_BUF_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R1_INV_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R2_INV_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y26__R2_INV_1 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y26__R3_BUF_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y27__R0_BUF_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R0_INV_0 (.A(tie_lo_T33Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y27__R1_BUF_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R1_INV_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R2_INV_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y27__R2_INV_1 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y27__R3_BUF_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y28__R0_BUF_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R0_INV_0 (.A(tie_lo_T33Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y28__R1_BUF_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R1_INV_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R2_INV_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y28__R2_INV_1 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y28__R3_BUF_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y29__R0_BUF_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R0_INV_0 (.A(tie_lo_T33Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y29__R1_BUF_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R1_INV_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R2_INV_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y29__R2_INV_1 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y29__R3_BUF_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y2__R0_BUF_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R0_INV_0 (.A(tie_lo_T33Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y2__R1_BUF_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R1_INV_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R2_INV_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y2__R2_INV_1 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y2__R3_BUF_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y30__R0_BUF_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R0_INV_0 (.A(tie_lo_T33Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y30__R1_BUF_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R1_INV_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R2_INV_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y30__R2_INV_1 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y30__R3_BUF_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y31__R0_BUF_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R0_INV_0 (.A(tie_lo_T33Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y31__R1_BUF_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R1_INV_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R2_INV_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y31__R2_INV_1 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y31__R3_BUF_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y32__R0_BUF_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R0_INV_0 (.A(tie_lo_T33Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y32__R1_BUF_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R1_INV_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R2_INV_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y32__R2_INV_1 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y32__R3_BUF_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y33__R0_BUF_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R0_INV_0 (.A(tie_lo_T33Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y33__R1_BUF_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R1_INV_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R2_INV_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y33__R2_INV_1 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y33__R3_BUF_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y34__R0_BUF_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R0_INV_0 (.A(tie_lo_T33Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y34__R1_BUF_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R1_INV_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R2_INV_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y34__R2_INV_1 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y34__R3_BUF_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y35__R0_BUF_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R0_INV_0 (.A(tie_lo_T33Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y35__R1_BUF_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R1_INV_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R2_INV_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y35__R2_INV_1 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y35__R3_BUF_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y36__R0_BUF_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R0_INV_0 (.A(tie_lo_T33Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y36__R1_BUF_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R1_INV_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R2_INV_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y36__R2_INV_1 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y36__R3_BUF_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y37__R0_BUF_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R0_INV_0 (.A(tie_lo_T33Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y37__R1_BUF_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R1_INV_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R2_INV_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y37__R2_INV_1 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y37__R3_BUF_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y38__R0_BUF_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R0_INV_0 (.A(tie_lo_T33Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y38__R1_BUF_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R1_INV_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R2_INV_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y38__R2_INV_1 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y38__R3_BUF_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y39__R0_BUF_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R0_INV_0 (.A(tie_lo_T33Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y39__R1_BUF_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R1_INV_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R2_INV_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y39__R2_INV_1 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y39__R3_BUF_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y3__R0_BUF_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R0_INV_0 (.A(tie_lo_T33Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y3__R1_BUF_0 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R1_INV_0 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R2_INV_0 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y3__R2_INV_1 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y3__R3_BUF_0 (.A(tie_lo_T33Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y40__R0_BUF_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R0_INV_0 (.A(tie_lo_T33Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y40__R1_BUF_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R1_INV_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R2_INV_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y40__R2_INV_1 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y40__R3_BUF_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y41__R0_BUF_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R0_INV_0 (.A(tie_lo_T33Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y41__R1_BUF_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R1_INV_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R2_INV_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y41__R2_INV_1 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y41__R3_BUF_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y42__R0_BUF_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R0_INV_0 (.A(tie_lo_T33Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y42__R1_BUF_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R1_INV_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R2_INV_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y42__R2_INV_1 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y42__R3_BUF_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y43__R0_BUF_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R0_INV_0 (.A(tie_lo_T33Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y43__R1_BUF_0 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R1_INV_0 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R2_INV_0 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y43__R2_INV_1 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y43__R3_BUF_0 (.A(tie_lo_T33Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y44__R0_BUF_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R0_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y44__R1_BUF_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R1_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R2_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y44__R2_INV_1 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y44__R3_BUF_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y45__R0_BUF_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R0_INV_0 (.A(tie_lo_T33Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y45__R1_BUF_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R1_INV_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R2_INV_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y45__R2_INV_1 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y45__R3_BUF_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y46__R0_BUF_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R0_INV_0 (.A(tie_lo_T33Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y46__R1_BUF_0 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R1_INV_0 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R2_INV_0 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y46__R2_INV_1 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y46__R3_BUF_0 (.A(tie_lo_T33Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y47__R0_BUF_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R0_INV_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y47__R1_BUF_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R1_INV_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R2_INV_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y47__R2_INV_1 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y47__R3_BUF_0 (.A(tie_lo_T33Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y48__R0_BUF_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R0_INV_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y48__R1_BUF_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R1_INV_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R2_INV_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y48__R2_INV_1 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y48__R3_BUF_0 (.A(tie_lo_T33Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y49__R0_BUF_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R0_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y49__R1_BUF_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R1_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R2_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y49__R2_INV_1 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y49__R3_BUF_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y4__R0_BUF_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R0_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y4__R1_BUF_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R1_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R2_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y4__R2_INV_1 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y4__R3_BUF_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y50__R0_BUF_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R0_INV_0 (.A(tie_lo_T33Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y50__R1_BUF_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R1_INV_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R2_INV_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y50__R2_INV_1 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y50__R3_BUF_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y51__R0_BUF_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R0_INV_0 (.A(tie_lo_T33Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y51__R1_BUF_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R1_INV_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R2_INV_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y51__R2_INV_1 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y51__R3_BUF_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y52__R0_BUF_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R0_INV_0 (.A(tie_lo_T33Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y52__R1_BUF_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R1_INV_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R2_INV_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y52__R2_INV_1 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y52__R3_BUF_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y53__R0_BUF_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R0_INV_0 (.A(tie_lo_T33Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y53__R1_BUF_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R1_INV_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R2_INV_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y53__R2_INV_1 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y53__R3_BUF_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y54__R0_BUF_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R0_INV_0 (.A(tie_lo_T33Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y54__R1_BUF_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R1_INV_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R2_INV_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y54__R2_INV_1 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y54__R3_BUF_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y55__R0_BUF_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R0_INV_0 (.A(tie_lo_T33Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y55__R1_BUF_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R1_INV_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R2_INV_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y55__R2_INV_1 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y55__R3_BUF_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y56__R0_BUF_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R0_INV_0 (.A(tie_lo_T33Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y56__R1_BUF_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R1_INV_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R2_INV_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y56__R2_INV_1 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y56__R3_BUF_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y57__R0_BUF_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R0_INV_0 (.A(tie_lo_T33Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y57__R1_BUF_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R1_INV_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R2_INV_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y57__R2_INV_1 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y57__R3_BUF_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y58__R0_BUF_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R0_INV_0 (.A(tie_lo_T33Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y58__R1_BUF_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R1_INV_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R2_INV_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y58__R2_INV_1 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y58__R3_BUF_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y59__R0_BUF_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R0_INV_0 (.A(tie_lo_T33Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y59__R1_BUF_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R1_INV_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R2_INV_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y59__R2_INV_1 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y59__R3_BUF_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y5__R0_BUF_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R0_INV_0 (.A(tie_lo_T33Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y5__R1_BUF_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R1_INV_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R2_INV_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y5__R2_INV_1 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y5__R3_BUF_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y60__R0_BUF_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R0_INV_0 (.A(tie_lo_T33Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y60__R1_BUF_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R1_INV_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R2_INV_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y60__R2_INV_1 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y60__R3_BUF_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y61__R0_BUF_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R0_INV_0 (.A(tie_lo_T33Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y61__R1_BUF_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R1_INV_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R2_INV_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y61__R2_INV_1 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y61__R3_BUF_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y62__R0_BUF_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R0_INV_0 (.A(tie_lo_T33Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y62__R1_BUF_0 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R1_INV_0 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R2_INV_0 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y62__R2_INV_1 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y62__R3_BUF_0 (.A(tie_lo_T33Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y63__R0_BUF_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R0_INV_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y63__R1_BUF_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R1_INV_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R2_INV_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y63__R2_INV_1 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y63__R3_BUF_0 (.A(tie_lo_T33Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y64__R0_BUF_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R0_INV_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y64__R1_BUF_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R1_INV_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R2_INV_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y64__R2_INV_1 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y64__R3_BUF_0 (.A(tie_lo_T33Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y65__R0_BUF_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R0_INV_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y65__R1_BUF_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R1_INV_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R2_INV_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y65__R2_INV_1 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y65__R3_BUF_0 (.A(tie_lo_T33Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y66__R0_BUF_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R0_INV_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y66__R1_BUF_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R1_INV_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R2_INV_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y66__R2_INV_1 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y66__R3_BUF_0 (.A(tie_lo_T33Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y67__R0_BUF_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R0_INV_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y67__R1_BUF_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R1_INV_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R2_INV_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y67__R2_INV_1 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y67__R3_BUF_0 (.A(tie_lo_T33Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y68__R0_BUF_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R0_INV_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y68__R1_BUF_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R1_INV_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R2_INV_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y68__R2_INV_1 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y68__R3_BUF_0 (.A(tie_lo_T33Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y69__R0_BUF_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R0_INV_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y69__R1_BUF_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R1_INV_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R2_INV_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y69__R2_INV_1 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y69__R3_BUF_0 (.A(tie_lo_T33Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y6__R0_BUF_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R0_INV_0 (.A(tie_lo_T33Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y6__R1_BUF_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R1_INV_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R2_INV_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y6__R2_INV_1 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y6__R3_BUF_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y70__R0_BUF_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R0_INV_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y70__R1_BUF_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R1_INV_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R2_INV_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y70__R2_INV_1 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y70__R3_BUF_0 (.A(tie_lo_T33Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y71__R0_BUF_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R0_INV_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y71__R1_BUF_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R1_INV_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R2_INV_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y71__R2_INV_1 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y71__R3_BUF_0 (.A(tie_lo_T33Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y72__R0_BUF_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R0_INV_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y72__R1_BUF_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R1_INV_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R2_INV_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y72__R2_INV_1 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y72__R3_BUF_0 (.A(tie_lo_T33Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y73__R0_BUF_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R0_INV_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y73__R1_BUF_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R1_INV_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R2_INV_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y73__R2_INV_1 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y73__R3_BUF_0 (.A(tie_lo_T33Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y74__R0_BUF_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R0_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y74__R1_BUF_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R1_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R2_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y74__R2_INV_1 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y74__R3_BUF_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y75__R0_BUF_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R0_INV_0 (.A(tie_lo_T33Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y75__R1_BUF_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R1_INV_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R2_INV_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y75__R2_INV_1 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y75__R3_BUF_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y76__R0_BUF_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R0_INV_0 (.A(tie_lo_T33Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y76__R1_BUF_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R1_INV_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R2_INV_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y76__R2_INV_1 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y76__R3_BUF_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y77__R0_BUF_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R0_INV_0 (.A(tie_lo_T33Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y77__R1_BUF_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R1_INV_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R2_INV_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y77__R2_INV_1 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y77__R3_BUF_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y78__R0_BUF_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R0_INV_0 (.A(tie_lo_T33Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y78__R1_BUF_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R1_INV_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R2_INV_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y78__R2_INV_1 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y78__R3_BUF_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y79__R0_BUF_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R0_INV_0 (.A(tie_lo_T33Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y79__R1_BUF_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R1_INV_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R2_INV_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y79__R2_INV_1 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y79__R3_BUF_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y7__R0_BUF_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R0_INV_0 (.A(tie_lo_T33Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y7__R1_BUF_0 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R1_INV_0 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R2_INV_0 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y7__R2_INV_1 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y7__R3_BUF_0 (.A(tie_lo_T33Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y80__R0_BUF_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R0_INV_0 (.A(tie_lo_T33Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y80__R1_BUF_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R1_INV_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R2_INV_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y80__R2_INV_1 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y80__R3_BUF_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y81__R0_BUF_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R0_INV_0 (.A(tie_lo_T33Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y81__R1_BUF_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R1_INV_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R2_INV_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y81__R2_INV_1 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y81__R3_BUF_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y82__R0_BUF_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R0_INV_0 (.A(tie_lo_T33Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y82__R1_BUF_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R1_INV_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R2_INV_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y82__R2_INV_1 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y82__R3_BUF_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y83__R0_BUF_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R0_INV_0 (.A(tie_lo_T33Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y83__R1_BUF_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R1_INV_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R2_INV_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y83__R2_INV_1 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y83__R3_BUF_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y84__R0_BUF_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R0_INV_0 (.A(tie_lo_T33Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y84__R1_BUF_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R1_INV_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R2_INV_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y84__R2_INV_1 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y84__R3_BUF_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y85__R0_BUF_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R0_INV_0 (.A(tie_lo_T33Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y85__R1_BUF_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R1_INV_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R2_INV_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y85__R2_INV_1 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y85__R3_BUF_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y86__R0_BUF_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R0_INV_0 (.A(tie_lo_T33Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y86__R1_BUF_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R1_INV_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R2_INV_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y86__R2_INV_1 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y86__R3_BUF_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y87__R0_BUF_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R0_INV_0 (.A(tie_lo_T33Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y87__R1_BUF_0 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R1_INV_0 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R2_INV_0 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y87__R2_INV_1 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y87__R3_BUF_0 (.A(tie_lo_T33Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y88__R0_BUF_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R0_INV_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y88__R1_BUF_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R1_INV_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R2_INV_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y88__R2_INV_1 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y88__R3_BUF_0 (.A(tie_lo_T33Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y89__R0_BUF_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R0_INV_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y89__R1_BUF_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R1_INV_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R2_INV_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y89__R2_INV_1 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y89__R3_BUF_0 (.A(tie_lo_T33Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y8__R0_BUF_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R0_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y8__R1_BUF_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R1_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R2_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y8__R2_INV_1 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y8__R3_BUF_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y9__R0_BUF_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R0_INV_0 (.A(tie_lo_T33Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y9__R1_BUF_0 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R1_INV_0 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T33Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R2_INV_0 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T33Y9__R2_INV_1 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T33Y9__R3_BUF_0 (.A(tie_lo_T33Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y0__R0_BUF_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R0_INV_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y0__R1_BUF_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R1_INV_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R2_INV_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y0__R2_INV_1 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y0__R3_BUF_0 (.A(tie_lo_T34Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y10__R0_BUF_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R0_INV_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y10__R1_BUF_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R1_INV_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R2_INV_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y10__R2_INV_1 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y10__R3_BUF_0 (.A(tie_lo_T34Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y11__R0_BUF_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R0_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y11__R1_BUF_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R1_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R2_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y11__R2_INV_1 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y11__R3_BUF_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y12__R0_BUF_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R0_INV_0 (.A(tie_lo_T34Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y12__R1_BUF_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R1_INV_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R2_INV_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y12__R2_INV_1 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y12__R3_BUF_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y13__R0_BUF_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R0_INV_0 (.A(tie_lo_T34Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y13__R1_BUF_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R1_INV_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R2_INV_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y13__R2_INV_1 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y13__R3_BUF_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y14__R0_BUF_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R0_INV_0 (.A(tie_lo_T34Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y14__R1_BUF_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R1_INV_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R2_INV_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y14__R2_INV_1 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y14__R3_BUF_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y15__R0_BUF_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R0_INV_0 (.A(tie_lo_T34Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y15__R1_BUF_0 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R1_INV_0 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R2_INV_0 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y15__R2_INV_1 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y15__R3_BUF_0 (.A(tie_lo_T34Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y16__R0_BUF_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R0_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y16__R1_BUF_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R1_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R2_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y16__R2_INV_1 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y16__R3_BUF_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y17__R0_BUF_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R0_INV_0 (.A(tie_lo_T34Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y17__R1_BUF_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R1_INV_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R2_INV_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y17__R2_INV_1 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y17__R3_BUF_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y18__R0_BUF_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R0_INV_0 (.A(tie_lo_T34Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y18__R1_BUF_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R1_INV_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R2_INV_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y18__R2_INV_1 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y18__R3_BUF_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y19__R0_BUF_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R0_INV_0 (.A(tie_lo_T34Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y19__R1_BUF_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R1_INV_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R2_INV_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y19__R2_INV_1 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y19__R3_BUF_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y1__R0_BUF_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R0_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y1__R1_BUF_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R1_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R2_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y1__R2_INV_1 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y1__R3_BUF_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y20__R0_BUF_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R0_INV_0 (.A(tie_lo_T34Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y20__R1_BUF_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R1_INV_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R2_INV_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y20__R2_INV_1 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y20__R3_BUF_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y21__R0_BUF_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R0_INV_0 (.A(tie_lo_T34Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y21__R1_BUF_0 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R1_INV_0 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R2_INV_0 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y21__R2_INV_1 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y21__R3_BUF_0 (.A(tie_lo_T34Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y22__R0_BUF_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R0_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y22__R1_BUF_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R1_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R2_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y22__R2_INV_1 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y22__R3_BUF_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y23__R0_BUF_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R0_INV_0 (.A(tie_lo_T34Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y23__R1_BUF_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R1_INV_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R2_INV_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y23__R2_INV_1 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y23__R3_BUF_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y24__R0_BUF_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R0_INV_0 (.A(tie_lo_T34Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y24__R1_BUF_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R1_INV_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R2_INV_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y24__R2_INV_1 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y24__R3_BUF_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y25__R0_BUF_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R0_INV_0 (.A(tie_lo_T34Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y25__R1_BUF_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R1_INV_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R2_INV_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y25__R2_INV_1 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y25__R3_BUF_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y26__R0_BUF_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R0_INV_0 (.A(tie_lo_T34Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y26__R1_BUF_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R1_INV_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R2_INV_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y26__R2_INV_1 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y26__R3_BUF_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y27__R0_BUF_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R0_INV_0 (.A(tie_lo_T34Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y27__R1_BUF_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R1_INV_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R2_INV_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y27__R2_INV_1 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y27__R3_BUF_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y28__R0_BUF_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R0_INV_0 (.A(tie_lo_T34Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y28__R1_BUF_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R1_INV_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R2_INV_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y28__R2_INV_1 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y28__R3_BUF_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y29__R0_BUF_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R0_INV_0 (.A(tie_lo_T34Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y29__R1_BUF_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R1_INV_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R2_INV_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y29__R2_INV_1 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y29__R3_BUF_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y2__R0_BUF_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R0_INV_0 (.A(tie_lo_T34Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y2__R1_BUF_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R1_INV_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R2_INV_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y2__R2_INV_1 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y2__R3_BUF_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y30__R0_BUF_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R0_INV_0 (.A(tie_lo_T34Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y30__R1_BUF_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R1_INV_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R2_INV_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y30__R2_INV_1 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y30__R3_BUF_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y31__R0_BUF_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R0_INV_0 (.A(tie_lo_T34Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y31__R1_BUF_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R1_INV_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R2_INV_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y31__R2_INV_1 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y31__R3_BUF_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y32__R0_BUF_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R0_INV_0 (.A(tie_lo_T34Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y32__R1_BUF_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R1_INV_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R2_INV_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y32__R2_INV_1 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y32__R3_BUF_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y33__R0_BUF_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R0_INV_0 (.A(tie_lo_T34Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y33__R1_BUF_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R1_INV_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R2_INV_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y33__R2_INV_1 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y33__R3_BUF_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y34__R0_BUF_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R0_INV_0 (.A(tie_lo_T34Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y34__R1_BUF_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R1_INV_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R2_INV_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y34__R2_INV_1 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y34__R3_BUF_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y35__R0_BUF_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R0_INV_0 (.A(tie_lo_T34Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y35__R1_BUF_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R1_INV_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R2_INV_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y35__R2_INV_1 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y35__R3_BUF_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y36__R0_BUF_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R0_INV_0 (.A(tie_lo_T34Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y36__R1_BUF_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R1_INV_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R2_INV_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y36__R2_INV_1 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y36__R3_BUF_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y37__R0_BUF_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R0_INV_0 (.A(tie_lo_T34Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y37__R1_BUF_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R1_INV_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R2_INV_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y37__R2_INV_1 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y37__R3_BUF_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y38__R0_BUF_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R0_INV_0 (.A(tie_lo_T34Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y38__R1_BUF_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R1_INV_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R2_INV_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y38__R2_INV_1 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y38__R3_BUF_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y39__R0_BUF_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R0_INV_0 (.A(tie_lo_T34Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y39__R1_BUF_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R1_INV_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R2_INV_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y39__R2_INV_1 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y39__R3_BUF_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y3__R0_BUF_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R0_INV_0 (.A(tie_lo_T34Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y3__R1_BUF_0 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R1_INV_0 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R2_INV_0 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y3__R2_INV_1 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y3__R3_BUF_0 (.A(tie_lo_T34Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y40__R0_BUF_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R0_INV_0 (.A(tie_lo_T34Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y40__R1_BUF_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R1_INV_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R2_INV_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y40__R2_INV_1 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y40__R3_BUF_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y41__R0_BUF_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R0_INV_0 (.A(tie_lo_T34Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y41__R1_BUF_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R1_INV_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R2_INV_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y41__R2_INV_1 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y41__R3_BUF_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y42__R0_BUF_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R0_INV_0 (.A(tie_lo_T34Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y42__R1_BUF_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R1_INV_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R2_INV_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y42__R2_INV_1 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y42__R3_BUF_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y43__R0_BUF_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R0_INV_0 (.A(tie_lo_T34Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y43__R1_BUF_0 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R1_INV_0 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R2_INV_0 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y43__R2_INV_1 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y43__R3_BUF_0 (.A(tie_lo_T34Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y44__R0_BUF_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R0_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y44__R1_BUF_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R1_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R2_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y44__R2_INV_1 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y44__R3_BUF_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y45__R0_BUF_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R0_INV_0 (.A(tie_lo_T34Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y45__R1_BUF_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R1_INV_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R2_INV_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y45__R2_INV_1 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y45__R3_BUF_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y46__R0_BUF_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R0_INV_0 (.A(tie_lo_T34Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y46__R1_BUF_0 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R1_INV_0 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R2_INV_0 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y46__R2_INV_1 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y46__R3_BUF_0 (.A(tie_lo_T34Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y47__R0_BUF_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R0_INV_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y47__R1_BUF_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R1_INV_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R2_INV_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y47__R2_INV_1 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y47__R3_BUF_0 (.A(tie_lo_T34Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y48__R0_BUF_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R0_INV_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y48__R1_BUF_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R1_INV_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R2_INV_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y48__R2_INV_1 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y48__R3_BUF_0 (.A(tie_lo_T34Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y49__R0_BUF_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R0_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y49__R1_BUF_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R1_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R2_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y49__R2_INV_1 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y49__R3_BUF_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y4__R0_BUF_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R0_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y4__R1_BUF_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R1_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R2_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y4__R2_INV_1 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y4__R3_BUF_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y50__R0_BUF_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R0_INV_0 (.A(tie_lo_T34Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y50__R1_BUF_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R1_INV_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R2_INV_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y50__R2_INV_1 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y50__R3_BUF_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y51__R0_BUF_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R0_INV_0 (.A(tie_lo_T34Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y51__R1_BUF_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R1_INV_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R2_INV_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y51__R2_INV_1 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y51__R3_BUF_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y52__R0_BUF_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R0_INV_0 (.A(tie_lo_T34Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y52__R1_BUF_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R1_INV_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R2_INV_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y52__R2_INV_1 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y52__R3_BUF_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y53__R0_BUF_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R0_INV_0 (.A(tie_lo_T34Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y53__R1_BUF_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R1_INV_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R2_INV_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y53__R2_INV_1 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y53__R3_BUF_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y54__R0_BUF_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R0_INV_0 (.A(tie_lo_T34Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y54__R1_BUF_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R1_INV_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R2_INV_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y54__R2_INV_1 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y54__R3_BUF_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y55__R0_BUF_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R0_INV_0 (.A(tie_lo_T34Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y55__R1_BUF_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R1_INV_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R2_INV_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y55__R2_INV_1 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y55__R3_BUF_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y56__R0_BUF_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R0_INV_0 (.A(tie_lo_T34Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y56__R1_BUF_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R1_INV_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R2_INV_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y56__R2_INV_1 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y56__R3_BUF_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y57__R0_BUF_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R0_INV_0 (.A(tie_lo_T34Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y57__R1_BUF_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R1_INV_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R2_INV_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y57__R2_INV_1 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y57__R3_BUF_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y58__R0_BUF_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R0_INV_0 (.A(tie_lo_T34Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y58__R1_BUF_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R1_INV_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R2_INV_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y58__R2_INV_1 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y58__R3_BUF_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y59__R0_BUF_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R0_INV_0 (.A(tie_lo_T34Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y59__R1_BUF_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R1_INV_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R2_INV_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y59__R2_INV_1 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y59__R3_BUF_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y5__R0_BUF_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R0_INV_0 (.A(tie_lo_T34Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y5__R1_BUF_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R1_INV_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R2_INV_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y5__R2_INV_1 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y5__R3_BUF_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y60__R0_BUF_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R0_INV_0 (.A(tie_lo_T34Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y60__R1_BUF_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R1_INV_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R2_INV_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y60__R2_INV_1 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y60__R3_BUF_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y61__R0_BUF_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R0_INV_0 (.A(tie_lo_T34Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y61__R1_BUF_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R1_INV_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R2_INV_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y61__R2_INV_1 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y61__R3_BUF_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y62__R0_BUF_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R0_INV_0 (.A(tie_lo_T34Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y62__R1_BUF_0 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R1_INV_0 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R2_INV_0 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y62__R2_INV_1 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y62__R3_BUF_0 (.A(tie_lo_T34Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y63__R0_BUF_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R0_INV_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y63__R1_BUF_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R1_INV_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R2_INV_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y63__R2_INV_1 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y63__R3_BUF_0 (.A(tie_lo_T34Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y64__R0_BUF_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R0_INV_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y64__R1_BUF_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R1_INV_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R2_INV_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y64__R2_INV_1 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y64__R3_BUF_0 (.A(tie_lo_T34Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y65__R0_BUF_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R0_INV_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y65__R1_BUF_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R1_INV_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R2_INV_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y65__R2_INV_1 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y65__R3_BUF_0 (.A(tie_lo_T34Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y66__R0_BUF_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R0_INV_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y66__R1_BUF_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R1_INV_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R2_INV_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y66__R2_INV_1 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y66__R3_BUF_0 (.A(tie_lo_T34Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y67__R0_BUF_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R0_INV_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y67__R1_BUF_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R1_INV_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R2_INV_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y67__R2_INV_1 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y67__R3_BUF_0 (.A(tie_lo_T34Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y68__R0_BUF_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R0_INV_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y68__R1_BUF_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R1_INV_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R2_INV_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y68__R2_INV_1 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y68__R3_BUF_0 (.A(tie_lo_T34Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y69__R0_BUF_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R0_INV_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y69__R1_BUF_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R1_INV_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R2_INV_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y69__R2_INV_1 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y69__R3_BUF_0 (.A(tie_lo_T34Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y6__R0_BUF_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R0_INV_0 (.A(tie_lo_T34Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y6__R1_BUF_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R1_INV_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R2_INV_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y6__R2_INV_1 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y6__R3_BUF_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y70__R0_BUF_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R0_INV_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y70__R1_BUF_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R1_INV_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R2_INV_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y70__R2_INV_1 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y70__R3_BUF_0 (.A(tie_lo_T34Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y71__R0_BUF_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R0_INV_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y71__R1_BUF_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R1_INV_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R2_INV_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y71__R2_INV_1 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y71__R3_BUF_0 (.A(tie_lo_T34Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y72__R0_BUF_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R0_INV_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y72__R1_BUF_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R1_INV_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R2_INV_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y72__R2_INV_1 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y72__R3_BUF_0 (.A(tie_lo_T34Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y73__R0_BUF_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R0_INV_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y73__R1_BUF_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R1_INV_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R2_INV_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y73__R2_INV_1 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y73__R3_BUF_0 (.A(tie_lo_T34Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y74__R0_BUF_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R0_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y74__R1_BUF_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R1_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R2_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y74__R2_INV_1 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y74__R3_BUF_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y75__R0_BUF_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R0_INV_0 (.A(tie_lo_T34Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y75__R1_BUF_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R1_INV_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R2_INV_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y75__R2_INV_1 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y75__R3_BUF_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y76__R0_BUF_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R0_INV_0 (.A(tie_lo_T34Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y76__R1_BUF_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R1_INV_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R2_INV_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y76__R2_INV_1 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y76__R3_BUF_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y77__R0_BUF_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R0_INV_0 (.A(tie_lo_T34Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y77__R1_BUF_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R1_INV_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R2_INV_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y77__R2_INV_1 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y77__R3_BUF_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y78__R0_BUF_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R0_INV_0 (.A(tie_lo_T34Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y78__R1_BUF_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R1_INV_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R2_INV_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y78__R2_INV_1 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y78__R3_BUF_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y79__R0_BUF_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R0_INV_0 (.A(tie_lo_T34Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y79__R1_BUF_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R1_INV_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R2_INV_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y79__R2_INV_1 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y79__R3_BUF_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y7__R0_BUF_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R0_INV_0 (.A(tie_lo_T34Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y7__R1_BUF_0 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R1_INV_0 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R2_INV_0 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y7__R2_INV_1 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y7__R3_BUF_0 (.A(tie_lo_T34Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y80__R0_BUF_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R0_INV_0 (.A(tie_lo_T34Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y80__R1_BUF_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R1_INV_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R2_INV_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y80__R2_INV_1 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y80__R3_BUF_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y81__R0_BUF_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R0_INV_0 (.A(tie_lo_T34Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y81__R1_BUF_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R1_INV_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R2_INV_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y81__R2_INV_1 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y81__R3_BUF_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y82__R0_BUF_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R0_INV_0 (.A(tie_lo_T34Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y82__R1_BUF_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R1_INV_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R2_INV_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y82__R2_INV_1 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y82__R3_BUF_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y83__R0_BUF_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R0_INV_0 (.A(tie_lo_T34Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y83__R1_BUF_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R1_INV_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R2_INV_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y83__R2_INV_1 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y83__R3_BUF_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y84__R0_BUF_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R0_INV_0 (.A(tie_lo_T34Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y84__R1_BUF_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R1_INV_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R2_INV_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y84__R2_INV_1 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y84__R3_BUF_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y85__R0_BUF_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R0_INV_0 (.A(tie_lo_T34Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y85__R1_BUF_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R1_INV_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R2_INV_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y85__R2_INV_1 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y85__R3_BUF_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y86__R0_BUF_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R0_INV_0 (.A(tie_lo_T34Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y86__R1_BUF_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R1_INV_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R2_INV_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y86__R2_INV_1 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y86__R3_BUF_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y87__R0_BUF_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R0_INV_0 (.A(tie_lo_T34Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y87__R1_BUF_0 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R1_INV_0 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R2_INV_0 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y87__R2_INV_1 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y87__R3_BUF_0 (.A(tie_lo_T34Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y88__R0_BUF_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R0_INV_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y88__R1_BUF_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R1_INV_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R2_INV_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y88__R2_INV_1 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y88__R3_BUF_0 (.A(tie_lo_T34Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y89__R0_BUF_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R0_INV_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y89__R1_BUF_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R1_INV_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R2_INV_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y89__R2_INV_1 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y89__R3_BUF_0 (.A(tie_lo_T34Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y8__R0_BUF_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R0_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y8__R1_BUF_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R1_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R2_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y8__R2_INV_1 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y8__R3_BUF_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y9__R0_BUF_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R0_INV_0 (.A(tie_lo_T34Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y9__R1_BUF_0 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R1_INV_0 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T34Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R2_INV_0 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T34Y9__R2_INV_1 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T34Y9__R3_BUF_0 (.A(tie_lo_T34Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y0__R0_BUF_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R0_INV_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y0__R1_BUF_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R1_INV_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R2_INV_0 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y0__R2_INV_1 (.A(tie_lo_T35Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y0__R3_BUF_0 (.A(clk), .X(clk_buf_T35Y0__R3_BUF_0_out));
  sky130_fd_sc_hd__clkbuf_4 T35Y10__R0_BUF_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R0_INV_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y10__R1_BUF_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R1_INV_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R2_INV_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y10__R2_INV_1 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y10__R3_BUF_0 (.A(tie_lo_T35Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y11__R0_BUF_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R0_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y11__R1_BUF_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R1_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R2_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y11__R2_INV_1 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y11__R3_BUF_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y12__R0_BUF_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R0_INV_0 (.A(tie_lo_T35Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y12__R1_BUF_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R1_INV_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R2_INV_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y12__R2_INV_1 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y12__R3_BUF_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y13__R0_BUF_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R0_INV_0 (.A(tie_lo_T35Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y13__R1_BUF_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R1_INV_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R2_INV_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y13__R2_INV_1 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y13__R3_BUF_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y14__R0_BUF_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R0_INV_0 (.A(tie_lo_T35Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y14__R1_BUF_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R1_INV_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R2_INV_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y14__R2_INV_1 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y14__R3_BUF_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y15__R0_BUF_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R0_INV_0 (.A(tie_lo_T35Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y15__R1_BUF_0 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R1_INV_0 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R2_INV_0 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y15__R2_INV_1 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y15__R3_BUF_0 (.A(tie_lo_T35Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y16__R0_BUF_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R0_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y16__R1_BUF_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R1_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R2_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y16__R2_INV_1 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y16__R3_BUF_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y17__R0_BUF_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R0_INV_0 (.A(tie_lo_T35Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y17__R1_BUF_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R1_INV_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R2_INV_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y17__R2_INV_1 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y17__R3_BUF_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y18__R0_BUF_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R0_INV_0 (.A(tie_lo_T35Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y18__R1_BUF_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R1_INV_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R2_INV_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y18__R2_INV_1 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y18__R3_BUF_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y19__R0_BUF_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R0_INV_0 (.A(tie_lo_T35Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y19__R1_BUF_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R1_INV_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R2_INV_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y19__R2_INV_1 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y19__R3_BUF_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y1__R0_BUF_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R0_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y1__R1_BUF_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R1_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R2_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y1__R2_INV_1 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y1__R3_BUF_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y20__R0_BUF_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R0_INV_0 (.A(tie_lo_T35Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y20__R1_BUF_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R1_INV_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R2_INV_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y20__R2_INV_1 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y20__R3_BUF_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y21__R0_BUF_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R0_INV_0 (.A(tie_lo_T35Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y21__R1_BUF_0 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R1_INV_0 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R2_INV_0 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y21__R2_INV_1 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y21__R3_BUF_0 (.A(tie_lo_T35Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y22__R0_BUF_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R0_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y22__R1_BUF_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R1_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R2_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y22__R2_INV_1 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y22__R3_BUF_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y23__R0_BUF_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R0_INV_0 (.A(tie_lo_T35Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y23__R1_BUF_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R1_INV_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R2_INV_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y23__R2_INV_1 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y23__R3_BUF_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y24__R0_BUF_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R0_INV_0 (.A(tie_lo_T35Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y24__R1_BUF_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R1_INV_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R2_INV_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y24__R2_INV_1 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y24__R3_BUF_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y25__R0_BUF_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R0_INV_0 (.A(tie_lo_T35Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y25__R1_BUF_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R1_INV_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R2_INV_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y25__R2_INV_1 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y25__R3_BUF_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y26__R0_BUF_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R0_INV_0 (.A(tie_lo_T35Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y26__R1_BUF_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R1_INV_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R2_INV_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y26__R2_INV_1 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y26__R3_BUF_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y27__R0_BUF_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R0_INV_0 (.A(tie_lo_T35Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y27__R1_BUF_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R1_INV_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R2_INV_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y27__R2_INV_1 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y27__R3_BUF_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y28__R0_BUF_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R0_INV_0 (.A(tie_lo_T35Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y28__R1_BUF_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R1_INV_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R2_INV_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y28__R2_INV_1 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y28__R3_BUF_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y29__R0_BUF_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R0_INV_0 (.A(tie_lo_T35Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y29__R1_BUF_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R1_INV_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R2_INV_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y29__R2_INV_1 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y29__R3_BUF_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y2__R0_BUF_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R0_INV_0 (.A(tie_lo_T35Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y2__R1_BUF_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R1_INV_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R2_INV_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y2__R2_INV_1 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y2__R3_BUF_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y30__R0_BUF_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R0_INV_0 (.A(tie_lo_T35Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y30__R1_BUF_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R1_INV_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R2_INV_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y30__R2_INV_1 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y30__R3_BUF_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y31__R0_BUF_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R0_INV_0 (.A(tie_lo_T35Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y31__R1_BUF_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R1_INV_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R2_INV_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y31__R2_INV_1 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y31__R3_BUF_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y32__R0_BUF_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R0_INV_0 (.A(tie_lo_T35Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y32__R1_BUF_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R1_INV_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R2_INV_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y32__R2_INV_1 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y32__R3_BUF_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y33__R0_BUF_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R0_INV_0 (.A(tie_lo_T35Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y33__R1_BUF_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R1_INV_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R2_INV_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y33__R2_INV_1 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y33__R3_BUF_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y34__R0_BUF_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R0_INV_0 (.A(tie_lo_T35Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y34__R1_BUF_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R1_INV_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R2_INV_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y34__R2_INV_1 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y34__R3_BUF_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y35__R0_BUF_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R0_INV_0 (.A(tie_lo_T35Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y35__R1_BUF_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R1_INV_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R2_INV_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y35__R2_INV_1 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y35__R3_BUF_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y36__R0_BUF_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R0_INV_0 (.A(tie_lo_T35Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y36__R1_BUF_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R1_INV_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R2_INV_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y36__R2_INV_1 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y36__R3_BUF_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y37__R0_BUF_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R0_INV_0 (.A(tie_lo_T35Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y37__R1_BUF_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R1_INV_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R2_INV_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y37__R2_INV_1 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y37__R3_BUF_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y38__R0_BUF_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R0_INV_0 (.A(tie_lo_T35Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y38__R1_BUF_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R1_INV_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R2_INV_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y38__R2_INV_1 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y38__R3_BUF_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y39__R0_BUF_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R0_INV_0 (.A(tie_lo_T35Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y39__R1_BUF_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R1_INV_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R2_INV_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y39__R2_INV_1 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y39__R3_BUF_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y3__R0_BUF_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R0_INV_0 (.A(tie_lo_T35Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y3__R1_BUF_0 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R1_INV_0 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R2_INV_0 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y3__R2_INV_1 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y3__R3_BUF_0 (.A(tie_lo_T35Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y40__R0_BUF_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R0_INV_0 (.A(tie_lo_T35Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y40__R1_BUF_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R1_INV_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R2_INV_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y40__R2_INV_1 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y40__R3_BUF_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y41__R0_BUF_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R0_INV_0 (.A(tie_lo_T35Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y41__R1_BUF_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R1_INV_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R2_INV_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y41__R2_INV_1 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y41__R3_BUF_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y42__R0_BUF_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R0_INV_0 (.A(tie_lo_T35Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y42__R1_BUF_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R1_INV_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R2_INV_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y42__R2_INV_1 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y42__R3_BUF_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y43__R0_BUF_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R0_INV_0 (.A(tie_lo_T35Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y43__R1_BUF_0 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R1_INV_0 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R2_INV_0 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y43__R2_INV_1 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y43__R3_BUF_0 (.A(tie_lo_T35Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y44__R0_BUF_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R0_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y44__R1_BUF_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R1_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R2_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y44__R2_INV_1 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y44__R3_BUF_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y45__R0_BUF_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R0_INV_0 (.A(tie_lo_T35Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y45__R1_BUF_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R1_INV_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R2_INV_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y45__R2_INV_1 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y45__R3_BUF_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y46__R0_BUF_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R0_INV_0 (.A(tie_lo_T35Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y46__R1_BUF_0 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R1_INV_0 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R2_INV_0 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y46__R2_INV_1 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y46__R3_BUF_0 (.A(tie_lo_T35Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y47__R0_BUF_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R0_INV_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y47__R1_BUF_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R1_INV_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R2_INV_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y47__R2_INV_1 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y47__R3_BUF_0 (.A(tie_lo_T35Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y48__R0_BUF_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R0_INV_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y48__R1_BUF_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R1_INV_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R2_INV_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y48__R2_INV_1 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y48__R3_BUF_0 (.A(tie_lo_T35Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y49__R0_BUF_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R0_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y49__R1_BUF_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R1_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R2_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y49__R2_INV_1 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y49__R3_BUF_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y4__R0_BUF_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R0_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y4__R1_BUF_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R1_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R2_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y4__R2_INV_1 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y4__R3_BUF_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y50__R0_BUF_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R0_INV_0 (.A(tie_lo_T35Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y50__R1_BUF_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R1_INV_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R2_INV_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y50__R2_INV_1 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y50__R3_BUF_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y51__R0_BUF_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R0_INV_0 (.A(tie_lo_T35Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y51__R1_BUF_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R1_INV_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R2_INV_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y51__R2_INV_1 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y51__R3_BUF_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y52__R0_BUF_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R0_INV_0 (.A(tie_lo_T35Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y52__R1_BUF_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R1_INV_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R2_INV_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y52__R2_INV_1 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y52__R3_BUF_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y53__R0_BUF_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R0_INV_0 (.A(tie_lo_T35Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y53__R1_BUF_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R1_INV_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R2_INV_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y53__R2_INV_1 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y53__R3_BUF_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y54__R0_BUF_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R0_INV_0 (.A(tie_lo_T35Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y54__R1_BUF_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R1_INV_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R2_INV_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y54__R2_INV_1 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y54__R3_BUF_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y55__R0_BUF_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R0_INV_0 (.A(tie_lo_T35Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y55__R1_BUF_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R1_INV_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R2_INV_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y55__R2_INV_1 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y55__R3_BUF_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y56__R0_BUF_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R0_INV_0 (.A(tie_lo_T35Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y56__R1_BUF_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R1_INV_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R2_INV_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y56__R2_INV_1 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y56__R3_BUF_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y57__R0_BUF_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R0_INV_0 (.A(tie_lo_T35Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y57__R1_BUF_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R1_INV_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R2_INV_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y57__R2_INV_1 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y57__R3_BUF_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y58__R0_BUF_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R0_INV_0 (.A(tie_lo_T35Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y58__R1_BUF_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R1_INV_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R2_INV_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y58__R2_INV_1 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y58__R3_BUF_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y59__R0_BUF_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R0_INV_0 (.A(tie_lo_T35Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y59__R1_BUF_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R1_INV_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R2_INV_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y59__R2_INV_1 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y59__R3_BUF_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y5__R0_BUF_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R0_INV_0 (.A(tie_lo_T35Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y5__R1_BUF_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R1_INV_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R2_INV_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y5__R2_INV_1 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y5__R3_BUF_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y60__R0_BUF_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R0_INV_0 (.A(tie_lo_T35Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y60__R1_BUF_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R1_INV_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R2_INV_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y60__R2_INV_1 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y60__R3_BUF_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y61__R0_BUF_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R0_INV_0 (.A(tie_lo_T35Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y61__R1_BUF_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R1_INV_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R2_INV_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y61__R2_INV_1 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y61__R3_BUF_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y62__R0_BUF_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R0_INV_0 (.A(tie_lo_T35Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y62__R1_BUF_0 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R1_INV_0 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R2_INV_0 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y62__R2_INV_1 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y62__R3_BUF_0 (.A(tie_lo_T35Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y63__R0_BUF_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R0_INV_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y63__R1_BUF_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R1_INV_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R2_INV_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y63__R2_INV_1 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y63__R3_BUF_0 (.A(tie_lo_T35Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y64__R0_BUF_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R0_INV_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y64__R1_BUF_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R1_INV_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R2_INV_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y64__R2_INV_1 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y64__R3_BUF_0 (.A(tie_lo_T35Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y65__R0_BUF_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R0_INV_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y65__R1_BUF_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R1_INV_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R2_INV_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y65__R2_INV_1 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y65__R3_BUF_0 (.A(tie_lo_T35Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y66__R0_BUF_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R0_INV_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y66__R1_BUF_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R1_INV_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R2_INV_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y66__R2_INV_1 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y66__R3_BUF_0 (.A(tie_lo_T35Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y67__R0_BUF_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R0_INV_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y67__R1_BUF_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R1_INV_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R2_INV_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y67__R2_INV_1 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y67__R3_BUF_0 (.A(tie_lo_T35Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y68__R0_BUF_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R0_INV_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y68__R1_BUF_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R1_INV_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R2_INV_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y68__R2_INV_1 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y68__R3_BUF_0 (.A(tie_lo_T35Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y69__R0_BUF_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R0_INV_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y69__R1_BUF_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R1_INV_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R2_INV_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y69__R2_INV_1 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y69__R3_BUF_0 (.A(tie_lo_T35Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y6__R0_BUF_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R0_INV_0 (.A(tie_lo_T35Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y6__R1_BUF_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R1_INV_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R2_INV_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y6__R2_INV_1 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y6__R3_BUF_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y70__R0_BUF_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R0_INV_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y70__R1_BUF_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R1_INV_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R2_INV_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y70__R2_INV_1 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y70__R3_BUF_0 (.A(tie_lo_T35Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y71__R0_BUF_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R0_INV_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y71__R1_BUF_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R1_INV_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R2_INV_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y71__R2_INV_1 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y71__R3_BUF_0 (.A(tie_lo_T35Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y72__R0_BUF_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R0_INV_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y72__R1_BUF_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R1_INV_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R2_INV_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y72__R2_INV_1 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y72__R3_BUF_0 (.A(tie_lo_T35Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y73__R0_BUF_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R0_INV_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y73__R1_BUF_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R1_INV_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R2_INV_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y73__R2_INV_1 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y73__R3_BUF_0 (.A(tie_lo_T35Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y74__R0_BUF_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R0_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y74__R1_BUF_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R1_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R2_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y74__R2_INV_1 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y74__R3_BUF_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y75__R0_BUF_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R0_INV_0 (.A(tie_lo_T35Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y75__R1_BUF_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R1_INV_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R2_INV_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y75__R2_INV_1 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y75__R3_BUF_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y76__R0_BUF_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R0_INV_0 (.A(tie_lo_T35Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y76__R1_BUF_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R1_INV_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R2_INV_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y76__R2_INV_1 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y76__R3_BUF_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y77__R0_BUF_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R0_INV_0 (.A(tie_lo_T35Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y77__R1_BUF_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R1_INV_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R2_INV_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y77__R2_INV_1 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y77__R3_BUF_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y78__R0_BUF_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R0_INV_0 (.A(tie_lo_T35Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y78__R1_BUF_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R1_INV_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R2_INV_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y78__R2_INV_1 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y78__R3_BUF_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y79__R0_BUF_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R0_INV_0 (.A(tie_lo_T35Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y79__R1_BUF_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R1_INV_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R2_INV_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y79__R2_INV_1 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y79__R3_BUF_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y7__R0_BUF_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R0_INV_0 (.A(tie_lo_T35Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y7__R1_BUF_0 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R1_INV_0 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R2_INV_0 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y7__R2_INV_1 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y7__R3_BUF_0 (.A(tie_lo_T35Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y80__R0_BUF_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R0_INV_0 (.A(tie_lo_T35Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y80__R1_BUF_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R1_INV_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R2_INV_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y80__R2_INV_1 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y80__R3_BUF_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y81__R0_BUF_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R0_INV_0 (.A(tie_lo_T35Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y81__R1_BUF_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R1_INV_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R2_INV_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y81__R2_INV_1 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y81__R3_BUF_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y82__R0_BUF_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R0_INV_0 (.A(tie_lo_T35Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y82__R1_BUF_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R1_INV_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R2_INV_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y82__R2_INV_1 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y82__R3_BUF_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y83__R0_BUF_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R0_INV_0 (.A(tie_lo_T35Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y83__R1_BUF_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R1_INV_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R2_INV_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y83__R2_INV_1 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y83__R3_BUF_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y84__R0_BUF_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R0_INV_0 (.A(tie_lo_T35Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y84__R1_BUF_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R1_INV_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R2_INV_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y84__R2_INV_1 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y84__R3_BUF_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y85__R0_BUF_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R0_INV_0 (.A(tie_lo_T35Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y85__R1_BUF_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R1_INV_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R2_INV_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y85__R2_INV_1 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y85__R3_BUF_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y86__R0_BUF_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R0_INV_0 (.A(tie_lo_T35Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y86__R1_BUF_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R1_INV_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R2_INV_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y86__R2_INV_1 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y86__R3_BUF_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y87__R0_BUF_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R0_INV_0 (.A(tie_lo_T35Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y87__R1_BUF_0 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R1_INV_0 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R2_INV_0 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y87__R2_INV_1 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y87__R3_BUF_0 (.A(tie_lo_T35Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y88__R0_BUF_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R0_INV_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y88__R1_BUF_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R1_INV_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R2_INV_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y88__R2_INV_1 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y88__R3_BUF_0 (.A(tie_lo_T35Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y89__R0_BUF_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R0_INV_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y89__R1_BUF_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R1_INV_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R2_INV_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y89__R2_INV_1 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y89__R3_BUF_0 (.A(tie_lo_T35Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y8__R0_BUF_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R0_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y8__R1_BUF_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R1_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R2_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y8__R2_INV_1 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y8__R3_BUF_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y9__R0_BUF_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R0_INV_0 (.A(tie_lo_T35Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y9__R1_BUF_0 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R1_INV_0 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T35Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R2_INV_0 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T35Y9__R2_INV_1 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T35Y9__R3_BUF_0 (.A(tie_lo_T35Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y0__R0_BUF_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R0_INV_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y0__R1_BUF_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R1_INV_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R2_INV_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y0__R2_INV_1 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y0__R3_BUF_0 (.A(tie_lo_T3Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y10__R0_BUF_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R0_INV_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y10__R1_BUF_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R1_INV_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R2_INV_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y10__R2_INV_1 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y10__R3_BUF_0 (.A(tie_lo_T3Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y11__R0_BUF_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R0_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y11__R1_BUF_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R1_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R2_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y11__R2_INV_1 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y11__R3_BUF_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y12__R0_BUF_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R0_INV_0 (.A(tie_lo_T3Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y12__R1_BUF_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R1_INV_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R2_INV_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y12__R2_INV_1 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y12__R3_BUF_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y13__R0_BUF_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R0_INV_0 (.A(tie_lo_T3Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y13__R1_BUF_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R1_INV_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R2_INV_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y13__R2_INV_1 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y13__R3_BUF_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y14__R0_BUF_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R0_INV_0 (.A(tie_lo_T3Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y14__R1_BUF_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R1_INV_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R2_INV_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y14__R2_INV_1 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y14__R3_BUF_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y15__R0_BUF_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R0_INV_0 (.A(tie_lo_T3Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y15__R1_BUF_0 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R1_INV_0 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R2_INV_0 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y15__R2_INV_1 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y15__R3_BUF_0 (.A(tie_lo_T3Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y16__R0_BUF_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R0_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y16__R1_BUF_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R1_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R2_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y16__R2_INV_1 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y16__R3_BUF_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y17__R0_BUF_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R0_INV_0 (.A(tie_lo_T3Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y17__R1_BUF_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R1_INV_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R2_INV_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y17__R2_INV_1 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y17__R3_BUF_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y18__R0_BUF_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R0_INV_0 (.A(tie_lo_T3Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y18__R1_BUF_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R1_INV_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R2_INV_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y18__R2_INV_1 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y18__R3_BUF_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y19__R0_BUF_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R0_INV_0 (.A(tie_lo_T3Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y19__R1_BUF_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R1_INV_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R2_INV_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y19__R2_INV_1 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y19__R3_BUF_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y1__R0_BUF_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R0_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y1__R1_BUF_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R1_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R2_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y1__R2_INV_1 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y1__R3_BUF_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y20__R0_BUF_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R0_INV_0 (.A(tie_lo_T3Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y20__R1_BUF_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R1_INV_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R2_INV_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y20__R2_INV_1 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y20__R3_BUF_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y21__R0_BUF_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R0_INV_0 (.A(tie_lo_T3Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y21__R1_BUF_0 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R1_INV_0 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R2_INV_0 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y21__R2_INV_1 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y21__R3_BUF_0 (.A(tie_lo_T3Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y22__R0_BUF_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R0_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y22__R1_BUF_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R1_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R2_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y22__R2_INV_1 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y22__R3_BUF_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y23__R0_BUF_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R0_INV_0 (.A(tie_lo_T3Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y23__R1_BUF_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R1_INV_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R2_INV_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y23__R2_INV_1 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y23__R3_BUF_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y24__R0_BUF_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R0_INV_0 (.A(tie_lo_T3Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y24__R1_BUF_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R1_INV_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R2_INV_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y24__R2_INV_1 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y24__R3_BUF_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y25__R0_BUF_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R0_INV_0 (.A(tie_lo_T3Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y25__R1_BUF_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R1_INV_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R2_INV_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y25__R2_INV_1 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y25__R3_BUF_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y26__R0_BUF_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R0_INV_0 (.A(tie_lo_T3Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y26__R1_BUF_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R1_INV_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R2_INV_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y26__R2_INV_1 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y26__R3_BUF_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y27__R0_BUF_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R0_INV_0 (.A(tie_lo_T3Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y27__R1_BUF_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R1_INV_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R2_INV_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y27__R2_INV_1 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y27__R3_BUF_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y28__R0_BUF_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R0_INV_0 (.A(tie_lo_T3Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y28__R1_BUF_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R1_INV_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R2_INV_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y28__R2_INV_1 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y28__R3_BUF_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y29__R0_BUF_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R0_INV_0 (.A(tie_lo_T3Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y29__R1_BUF_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R1_INV_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R2_INV_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y29__R2_INV_1 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y29__R3_BUF_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y2__R0_BUF_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R0_INV_0 (.A(tie_lo_T3Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y2__R1_BUF_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R1_INV_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R2_INV_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y2__R2_INV_1 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y2__R3_BUF_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y30__R0_BUF_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R0_INV_0 (.A(tie_lo_T3Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y30__R1_BUF_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R1_INV_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R2_INV_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y30__R2_INV_1 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y30__R3_BUF_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y31__R0_BUF_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R0_INV_0 (.A(tie_lo_T3Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y31__R1_BUF_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R1_INV_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R2_INV_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y31__R2_INV_1 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y31__R3_BUF_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y32__R0_BUF_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R0_INV_0 (.A(tie_lo_T3Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y32__R1_BUF_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R1_INV_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R2_INV_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y32__R2_INV_1 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y32__R3_BUF_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y33__R0_BUF_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R0_INV_0 (.A(tie_lo_T3Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y33__R1_BUF_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R1_INV_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R2_INV_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y33__R2_INV_1 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y33__R3_BUF_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y34__R0_BUF_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R0_INV_0 (.A(tie_lo_T3Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y34__R1_BUF_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R1_INV_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R2_INV_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y34__R2_INV_1 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y34__R3_BUF_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y35__R0_BUF_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R0_INV_0 (.A(tie_lo_T3Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y35__R1_BUF_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R1_INV_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R2_INV_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y35__R2_INV_1 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y35__R3_BUF_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y36__R0_BUF_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R0_INV_0 (.A(tie_lo_T3Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y36__R1_BUF_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R1_INV_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R2_INV_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y36__R2_INV_1 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y36__R3_BUF_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y37__R0_BUF_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R0_INV_0 (.A(tie_lo_T3Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y37__R1_BUF_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R1_INV_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R2_INV_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y37__R2_INV_1 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y37__R3_BUF_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y38__R0_BUF_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R0_INV_0 (.A(tie_lo_T3Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y38__R1_BUF_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R1_INV_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R2_INV_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y38__R2_INV_1 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y38__R3_BUF_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y39__R0_BUF_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R0_INV_0 (.A(tie_lo_T3Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y39__R1_BUF_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R1_INV_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R2_INV_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y39__R2_INV_1 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y39__R3_BUF_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y3__R0_BUF_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R0_INV_0 (.A(tie_lo_T3Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y3__R1_BUF_0 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R1_INV_0 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R2_INV_0 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y3__R2_INV_1 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y3__R3_BUF_0 (.A(tie_lo_T3Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y40__R0_BUF_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R0_INV_0 (.A(tie_lo_T3Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y40__R1_BUF_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R1_INV_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R2_INV_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y40__R2_INV_1 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y40__R3_BUF_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y41__R0_BUF_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R0_INV_0 (.A(tie_lo_T3Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y41__R1_BUF_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R1_INV_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R2_INV_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y41__R2_INV_1 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y41__R3_BUF_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y42__R0_BUF_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R0_INV_0 (.A(tie_lo_T3Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y42__R1_BUF_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R1_INV_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R2_INV_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y42__R2_INV_1 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y42__R3_BUF_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y43__R0_BUF_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R0_INV_0 (.A(tie_lo_T3Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y43__R1_BUF_0 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R1_INV_0 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R2_INV_0 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y43__R2_INV_1 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y43__R3_BUF_0 (.A(tie_lo_T3Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y44__R0_BUF_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R0_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y44__R1_BUF_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R1_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R2_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y44__R2_INV_1 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y44__R3_BUF_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y45__R0_BUF_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R0_INV_0 (.A(tie_lo_T3Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y45__R1_BUF_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R1_INV_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R2_INV_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y45__R2_INV_1 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y45__R3_BUF_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y46__R0_BUF_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R0_INV_0 (.A(tie_lo_T3Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y46__R1_BUF_0 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R1_INV_0 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R2_INV_0 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y46__R2_INV_1 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y46__R3_BUF_0 (.A(tie_lo_T3Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y47__R0_BUF_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R0_INV_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y47__R1_BUF_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R1_INV_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R2_INV_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y47__R2_INV_1 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y47__R3_BUF_0 (.A(tie_lo_T3Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y48__R0_BUF_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R0_INV_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y48__R1_BUF_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R1_INV_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R2_INV_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y48__R2_INV_1 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y48__R3_BUF_0 (.A(tie_lo_T3Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y49__R0_BUF_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R0_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y49__R1_BUF_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R1_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R2_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y49__R2_INV_1 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y49__R3_BUF_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y4__R0_BUF_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R0_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y4__R1_BUF_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R1_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R2_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y4__R2_INV_1 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y4__R3_BUF_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y50__R0_BUF_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R0_INV_0 (.A(tie_lo_T3Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y50__R1_BUF_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R1_INV_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R2_INV_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y50__R2_INV_1 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y50__R3_BUF_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y51__R0_BUF_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R0_INV_0 (.A(tie_lo_T3Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y51__R1_BUF_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R1_INV_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R2_INV_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y51__R2_INV_1 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y51__R3_BUF_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y52__R0_BUF_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R0_INV_0 (.A(tie_lo_T3Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y52__R1_BUF_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R1_INV_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R2_INV_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y52__R2_INV_1 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y52__R3_BUF_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y53__R0_BUF_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R0_INV_0 (.A(tie_lo_T3Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y53__R1_BUF_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R1_INV_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R2_INV_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y53__R2_INV_1 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y53__R3_BUF_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y54__R0_BUF_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R0_INV_0 (.A(tie_lo_T3Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y54__R1_BUF_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R1_INV_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R2_INV_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y54__R2_INV_1 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y54__R3_BUF_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y55__R0_BUF_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R0_INV_0 (.A(tie_lo_T3Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y55__R1_BUF_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R1_INV_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R2_INV_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y55__R2_INV_1 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y55__R3_BUF_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y56__R0_BUF_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R0_INV_0 (.A(tie_lo_T3Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y56__R1_BUF_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R1_INV_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R2_INV_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y56__R2_INV_1 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y56__R3_BUF_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y57__R0_BUF_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R0_INV_0 (.A(tie_lo_T3Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y57__R1_BUF_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R1_INV_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R2_INV_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y57__R2_INV_1 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y57__R3_BUF_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y58__R0_BUF_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R0_INV_0 (.A(tie_lo_T3Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y58__R1_BUF_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R1_INV_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R2_INV_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y58__R2_INV_1 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y58__R3_BUF_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y59__R0_BUF_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R0_INV_0 (.A(tie_lo_T3Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y59__R1_BUF_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R1_INV_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R2_INV_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y59__R2_INV_1 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y59__R3_BUF_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y5__R0_BUF_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R0_INV_0 (.A(tie_lo_T3Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y5__R1_BUF_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R1_INV_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R2_INV_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y5__R2_INV_1 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y5__R3_BUF_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y60__R0_BUF_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R0_INV_0 (.A(tie_lo_T3Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y60__R1_BUF_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R1_INV_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R2_INV_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y60__R2_INV_1 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y60__R3_BUF_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y61__R0_BUF_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R0_INV_0 (.A(tie_lo_T3Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y61__R1_BUF_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R1_INV_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R2_INV_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y61__R2_INV_1 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y61__R3_BUF_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y62__R0_BUF_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R0_INV_0 (.A(tie_lo_T3Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y62__R1_BUF_0 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R1_INV_0 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R2_INV_0 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y62__R2_INV_1 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y62__R3_BUF_0 (.A(tie_lo_T3Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y63__R0_BUF_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R0_INV_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y63__R1_BUF_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R1_INV_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R2_INV_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y63__R2_INV_1 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y63__R3_BUF_0 (.A(tie_lo_T3Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y64__R0_BUF_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R0_INV_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y64__R1_BUF_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R1_INV_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R2_INV_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y64__R2_INV_1 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y64__R3_BUF_0 (.A(tie_lo_T3Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y65__R0_BUF_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R0_INV_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y65__R1_BUF_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R1_INV_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R2_INV_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y65__R2_INV_1 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y65__R3_BUF_0 (.A(tie_lo_T3Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y66__R0_BUF_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R0_INV_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y66__R1_BUF_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R1_INV_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R2_INV_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y66__R2_INV_1 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y66__R3_BUF_0 (.A(tie_lo_T3Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y67__R0_BUF_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R0_INV_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y67__R1_BUF_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R1_INV_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R2_INV_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y67__R2_INV_1 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y67__R3_BUF_0 (.A(tie_lo_T3Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y68__R0_BUF_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R0_INV_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y68__R1_BUF_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R1_INV_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R2_INV_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y68__R2_INV_1 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y68__R3_BUF_0 (.A(tie_lo_T3Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y69__R0_BUF_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R0_INV_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y69__R1_BUF_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R1_INV_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R2_INV_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y69__R2_INV_1 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y69__R3_BUF_0 (.A(tie_lo_T3Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y6__R0_BUF_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R0_INV_0 (.A(tie_lo_T3Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y6__R1_BUF_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R1_INV_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R2_INV_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y6__R2_INV_1 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y6__R3_BUF_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y70__R0_BUF_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R0_INV_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y70__R1_BUF_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R1_INV_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R2_INV_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y70__R2_INV_1 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y70__R3_BUF_0 (.A(tie_lo_T3Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y71__R0_BUF_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R0_INV_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y71__R1_BUF_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R1_INV_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R2_INV_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y71__R2_INV_1 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y71__R3_BUF_0 (.A(tie_lo_T3Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y72__R0_BUF_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R0_INV_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y72__R1_BUF_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R1_INV_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R2_INV_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y72__R2_INV_1 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y72__R3_BUF_0 (.A(tie_lo_T3Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y73__R0_BUF_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R0_INV_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y73__R1_BUF_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R1_INV_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R2_INV_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y73__R2_INV_1 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y73__R3_BUF_0 (.A(tie_lo_T3Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y74__R0_BUF_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R0_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y74__R1_BUF_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R1_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R2_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y74__R2_INV_1 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y74__R3_BUF_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y75__R0_BUF_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R0_INV_0 (.A(tie_lo_T3Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y75__R1_BUF_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R1_INV_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R2_INV_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y75__R2_INV_1 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y75__R3_BUF_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y76__R0_BUF_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R0_INV_0 (.A(tie_lo_T3Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y76__R1_BUF_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R1_INV_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R2_INV_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y76__R2_INV_1 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y76__R3_BUF_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y77__R0_BUF_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R0_INV_0 (.A(tie_lo_T3Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y77__R1_BUF_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R1_INV_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R2_INV_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y77__R2_INV_1 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y77__R3_BUF_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y78__R0_BUF_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R0_INV_0 (.A(tie_lo_T3Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y78__R1_BUF_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R1_INV_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R2_INV_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y78__R2_INV_1 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y78__R3_BUF_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y79__R0_BUF_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R0_INV_0 (.A(tie_lo_T3Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y79__R1_BUF_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R1_INV_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R2_INV_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y79__R2_INV_1 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y79__R3_BUF_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y7__R0_BUF_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R0_INV_0 (.A(tie_lo_T3Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y7__R1_BUF_0 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R1_INV_0 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R2_INV_0 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y7__R2_INV_1 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y7__R3_BUF_0 (.A(tie_lo_T3Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y80__R0_BUF_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R0_INV_0 (.A(tie_lo_T3Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y80__R1_BUF_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R1_INV_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R2_INV_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y80__R2_INV_1 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y80__R3_BUF_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y81__R0_BUF_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R0_INV_0 (.A(tie_lo_T3Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y81__R1_BUF_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R1_INV_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R2_INV_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y81__R2_INV_1 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y81__R3_BUF_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y82__R0_BUF_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R0_INV_0 (.A(tie_lo_T3Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y82__R1_BUF_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R1_INV_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R2_INV_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y82__R2_INV_1 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y82__R3_BUF_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y83__R0_BUF_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R0_INV_0 (.A(tie_lo_T3Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y83__R1_BUF_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R1_INV_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R2_INV_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y83__R2_INV_1 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y83__R3_BUF_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y84__R0_BUF_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R0_INV_0 (.A(tie_lo_T3Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y84__R1_BUF_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R1_INV_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R2_INV_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y84__R2_INV_1 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y84__R3_BUF_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y85__R0_BUF_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R0_INV_0 (.A(tie_lo_T3Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y85__R1_BUF_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R1_INV_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R2_INV_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y85__R2_INV_1 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y85__R3_BUF_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y86__R0_BUF_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R0_INV_0 (.A(tie_lo_T3Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y86__R1_BUF_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R1_INV_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R2_INV_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y86__R2_INV_1 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y86__R3_BUF_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y87__R0_BUF_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R0_INV_0 (.A(tie_lo_T3Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y87__R1_BUF_0 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R1_INV_0 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R2_INV_0 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y87__R2_INV_1 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y87__R3_BUF_0 (.A(tie_lo_T3Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y88__R0_BUF_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R0_INV_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y88__R1_BUF_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R1_INV_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R2_INV_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y88__R2_INV_1 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y88__R3_BUF_0 (.A(tie_lo_T3Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y89__R0_BUF_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R0_INV_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y89__R1_BUF_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R1_INV_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R2_INV_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y89__R2_INV_1 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y89__R3_BUF_0 (.A(tie_lo_T3Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y8__R0_BUF_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R0_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y8__R1_BUF_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R1_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R2_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y8__R2_INV_1 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y8__R3_BUF_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y9__R0_BUF_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R0_INV_0 (.A(tie_lo_T3Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y9__R1_BUF_0 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R1_INV_0 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T3Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R2_INV_0 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T3Y9__R2_INV_1 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T3Y9__R3_BUF_0 (.A(tie_lo_T3Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y0__R0_BUF_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R0_INV_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y0__R1_BUF_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R1_INV_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R2_INV_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y0__R2_INV_1 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y0__R3_BUF_0 (.A(tie_lo_T4Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y10__R0_BUF_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R0_INV_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y10__R1_BUF_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R1_INV_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R2_INV_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y10__R2_INV_1 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y10__R3_BUF_0 (.A(tie_lo_T4Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y11__R0_BUF_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R0_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y11__R1_BUF_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R1_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R2_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y11__R2_INV_1 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y11__R3_BUF_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y12__R0_BUF_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R0_INV_0 (.A(tie_lo_T4Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y12__R1_BUF_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R1_INV_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R2_INV_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y12__R2_INV_1 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y12__R3_BUF_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y13__R0_BUF_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R0_INV_0 (.A(tie_lo_T4Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y13__R1_BUF_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R1_INV_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R2_INV_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y13__R2_INV_1 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y13__R3_BUF_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y14__R0_BUF_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R0_INV_0 (.A(tie_lo_T4Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y14__R1_BUF_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R1_INV_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R2_INV_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y14__R2_INV_1 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y14__R3_BUF_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y15__R0_BUF_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R0_INV_0 (.A(tie_lo_T4Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y15__R1_BUF_0 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R1_INV_0 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R2_INV_0 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y15__R2_INV_1 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y15__R3_BUF_0 (.A(tie_lo_T4Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y16__R0_BUF_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R0_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y16__R1_BUF_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R1_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R2_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y16__R2_INV_1 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y16__R3_BUF_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y17__R0_BUF_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R0_INV_0 (.A(tie_lo_T4Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y17__R1_BUF_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R1_INV_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R2_INV_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y17__R2_INV_1 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y17__R3_BUF_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y18__R0_BUF_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R0_INV_0 (.A(tie_lo_T4Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y18__R1_BUF_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R1_INV_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R2_INV_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y18__R2_INV_1 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y18__R3_BUF_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y19__R0_BUF_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R0_INV_0 (.A(tie_lo_T4Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y19__R1_BUF_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R1_INV_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R2_INV_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y19__R2_INV_1 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y19__R3_BUF_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y1__R0_BUF_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R0_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y1__R1_BUF_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R1_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R2_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y1__R2_INV_1 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y1__R3_BUF_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y20__R0_BUF_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R0_INV_0 (.A(tie_lo_T4Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y20__R1_BUF_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R1_INV_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R2_INV_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y20__R2_INV_1 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y20__R3_BUF_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y21__R0_BUF_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R0_INV_0 (.A(tie_lo_T4Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y21__R1_BUF_0 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R1_INV_0 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R2_INV_0 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y21__R2_INV_1 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y21__R3_BUF_0 (.A(tie_lo_T4Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y22__R0_BUF_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R0_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y22__R1_BUF_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R1_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R2_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y22__R2_INV_1 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y22__R3_BUF_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y23__R0_BUF_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R0_INV_0 (.A(tie_lo_T4Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y23__R1_BUF_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R1_INV_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R2_INV_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y23__R2_INV_1 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y23__R3_BUF_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y24__R0_BUF_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R0_INV_0 (.A(tie_lo_T4Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y24__R1_BUF_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R1_INV_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R2_INV_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y24__R2_INV_1 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y24__R3_BUF_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y25__R0_BUF_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R0_INV_0 (.A(tie_lo_T4Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y25__R1_BUF_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R1_INV_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R2_INV_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y25__R2_INV_1 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y25__R3_BUF_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y26__R0_BUF_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R0_INV_0 (.A(tie_lo_T4Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y26__R1_BUF_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R1_INV_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R2_INV_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y26__R2_INV_1 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y26__R3_BUF_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y27__R0_BUF_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R0_INV_0 (.A(tie_lo_T4Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y27__R1_BUF_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R1_INV_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R2_INV_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y27__R2_INV_1 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y27__R3_BUF_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y28__R0_BUF_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R0_INV_0 (.A(tie_lo_T4Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y28__R1_BUF_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R1_INV_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R2_INV_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y28__R2_INV_1 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y28__R3_BUF_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y29__R0_BUF_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R0_INV_0 (.A(tie_lo_T4Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y29__R1_BUF_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R1_INV_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R2_INV_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y29__R2_INV_1 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y29__R3_BUF_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y2__R0_BUF_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R0_INV_0 (.A(tie_lo_T4Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y2__R1_BUF_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R1_INV_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R2_INV_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y2__R2_INV_1 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y2__R3_BUF_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y30__R0_BUF_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R0_INV_0 (.A(tie_lo_T4Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y30__R1_BUF_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R1_INV_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R2_INV_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y30__R2_INV_1 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y30__R3_BUF_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y31__R0_BUF_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R0_INV_0 (.A(tie_lo_T4Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y31__R1_BUF_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R1_INV_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R2_INV_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y31__R2_INV_1 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y31__R3_BUF_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y32__R0_BUF_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R0_INV_0 (.A(tie_lo_T4Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y32__R1_BUF_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R1_INV_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R2_INV_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y32__R2_INV_1 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y32__R3_BUF_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y33__R0_BUF_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R0_INV_0 (.A(tie_lo_T4Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y33__R1_BUF_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R1_INV_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R2_INV_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y33__R2_INV_1 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y33__R3_BUF_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y34__R0_BUF_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R0_INV_0 (.A(tie_lo_T4Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y34__R1_BUF_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R1_INV_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R2_INV_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y34__R2_INV_1 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y34__R3_BUF_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y35__R0_BUF_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R0_INV_0 (.A(tie_lo_T4Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y35__R1_BUF_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R1_INV_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R2_INV_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y35__R2_INV_1 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y35__R3_BUF_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y36__R0_BUF_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R0_INV_0 (.A(tie_lo_T4Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y36__R1_BUF_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R1_INV_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R2_INV_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y36__R2_INV_1 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y36__R3_BUF_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y37__R0_BUF_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R0_INV_0 (.A(tie_lo_T4Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y37__R1_BUF_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R1_INV_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R2_INV_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y37__R2_INV_1 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y37__R3_BUF_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y38__R0_BUF_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R0_INV_0 (.A(tie_lo_T4Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y38__R1_BUF_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R1_INV_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R2_INV_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y38__R2_INV_1 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y38__R3_BUF_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y39__R0_BUF_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R0_INV_0 (.A(tie_lo_T4Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y39__R1_BUF_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R1_INV_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R2_INV_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y39__R2_INV_1 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y39__R3_BUF_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y3__R0_BUF_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R0_INV_0 (.A(tie_lo_T4Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y3__R1_BUF_0 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R1_INV_0 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R2_INV_0 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y3__R2_INV_1 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y3__R3_BUF_0 (.A(tie_lo_T4Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y40__R0_BUF_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R0_INV_0 (.A(tie_lo_T4Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y40__R1_BUF_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R1_INV_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R2_INV_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y40__R2_INV_1 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y40__R3_BUF_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y41__R0_BUF_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R0_INV_0 (.A(tie_lo_T4Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y41__R1_BUF_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R1_INV_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R2_INV_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y41__R2_INV_1 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y41__R3_BUF_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y42__R0_BUF_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R0_INV_0 (.A(tie_lo_T4Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y42__R1_BUF_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R1_INV_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R2_INV_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y42__R2_INV_1 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y42__R3_BUF_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y43__R0_BUF_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R0_INV_0 (.A(tie_lo_T4Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y43__R1_BUF_0 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R1_INV_0 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R2_INV_0 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y43__R2_INV_1 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y43__R3_BUF_0 (.A(tie_lo_T4Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y44__R0_BUF_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R0_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y44__R1_BUF_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R1_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R2_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y44__R2_INV_1 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y44__R3_BUF_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y45__R0_BUF_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R0_INV_0 (.A(tie_lo_T4Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y45__R1_BUF_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R1_INV_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R2_INV_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y45__R2_INV_1 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y45__R3_BUF_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y46__R0_BUF_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R0_INV_0 (.A(tie_lo_T4Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y46__R1_BUF_0 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R1_INV_0 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R2_INV_0 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y46__R2_INV_1 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y46__R3_BUF_0 (.A(tie_lo_T4Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y47__R0_BUF_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R0_INV_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y47__R1_BUF_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R1_INV_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R2_INV_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y47__R2_INV_1 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y47__R3_BUF_0 (.A(tie_lo_T4Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y48__R0_BUF_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R0_INV_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y48__R1_BUF_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R1_INV_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R2_INV_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y48__R2_INV_1 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y48__R3_BUF_0 (.A(tie_lo_T4Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y49__R0_BUF_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R0_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y49__R1_BUF_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R1_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R2_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y49__R2_INV_1 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y49__R3_BUF_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y4__R0_BUF_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R0_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y4__R1_BUF_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R1_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R2_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y4__R2_INV_1 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y4__R3_BUF_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y50__R0_BUF_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R0_INV_0 (.A(tie_lo_T4Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y50__R1_BUF_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R1_INV_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R2_INV_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y50__R2_INV_1 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y50__R3_BUF_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y51__R0_BUF_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R0_INV_0 (.A(tie_lo_T4Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y51__R1_BUF_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R1_INV_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R2_INV_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y51__R2_INV_1 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y51__R3_BUF_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y52__R0_BUF_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R0_INV_0 (.A(tie_lo_T4Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y52__R1_BUF_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R1_INV_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R2_INV_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y52__R2_INV_1 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y52__R3_BUF_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y53__R0_BUF_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R0_INV_0 (.A(tie_lo_T4Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y53__R1_BUF_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R1_INV_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R2_INV_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y53__R2_INV_1 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y53__R3_BUF_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y54__R0_BUF_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R0_INV_0 (.A(tie_lo_T4Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y54__R1_BUF_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R1_INV_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R2_INV_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y54__R2_INV_1 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y54__R3_BUF_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y55__R0_BUF_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R0_INV_0 (.A(tie_lo_T4Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y55__R1_BUF_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R1_INV_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R2_INV_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y55__R2_INV_1 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y55__R3_BUF_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y56__R0_BUF_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R0_INV_0 (.A(tie_lo_T4Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y56__R1_BUF_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R1_INV_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R2_INV_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y56__R2_INV_1 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y56__R3_BUF_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y57__R0_BUF_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R0_INV_0 (.A(tie_lo_T4Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y57__R1_BUF_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R1_INV_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R2_INV_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y57__R2_INV_1 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y57__R3_BUF_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y58__R0_BUF_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R0_INV_0 (.A(tie_lo_T4Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y58__R1_BUF_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R1_INV_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R2_INV_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y58__R2_INV_1 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y58__R3_BUF_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y59__R0_BUF_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R0_INV_0 (.A(tie_lo_T4Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y59__R1_BUF_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R1_INV_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R2_INV_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y59__R2_INV_1 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y59__R3_BUF_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y5__R0_BUF_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R0_INV_0 (.A(tie_lo_T4Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y5__R1_BUF_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R1_INV_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R2_INV_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y5__R2_INV_1 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y5__R3_BUF_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y60__R0_BUF_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R0_INV_0 (.A(tie_lo_T4Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y60__R1_BUF_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R1_INV_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R2_INV_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y60__R2_INV_1 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y60__R3_BUF_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y61__R0_BUF_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R0_INV_0 (.A(tie_lo_T4Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y61__R1_BUF_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R1_INV_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R2_INV_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y61__R2_INV_1 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y61__R3_BUF_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y62__R0_BUF_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R0_INV_0 (.A(tie_lo_T4Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y62__R1_BUF_0 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R1_INV_0 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R2_INV_0 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y62__R2_INV_1 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y62__R3_BUF_0 (.A(tie_lo_T4Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y63__R0_BUF_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R0_INV_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y63__R1_BUF_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R1_INV_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R2_INV_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y63__R2_INV_1 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y63__R3_BUF_0 (.A(tie_lo_T4Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y64__R0_BUF_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R0_INV_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y64__R1_BUF_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R1_INV_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R2_INV_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y64__R2_INV_1 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y64__R3_BUF_0 (.A(tie_lo_T4Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y65__R0_BUF_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R0_INV_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y65__R1_BUF_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R1_INV_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R2_INV_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y65__R2_INV_1 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y65__R3_BUF_0 (.A(tie_lo_T4Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y66__R0_BUF_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R0_INV_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y66__R1_BUF_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R1_INV_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R2_INV_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y66__R2_INV_1 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y66__R3_BUF_0 (.A(tie_lo_T4Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y67__R0_BUF_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R0_INV_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y67__R1_BUF_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R1_INV_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R2_INV_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y67__R2_INV_1 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y67__R3_BUF_0 (.A(tie_lo_T4Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y68__R0_BUF_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R0_INV_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y68__R1_BUF_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R1_INV_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R2_INV_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y68__R2_INV_1 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y68__R3_BUF_0 (.A(tie_lo_T4Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y69__R0_BUF_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R0_INV_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y69__R1_BUF_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R1_INV_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R2_INV_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y69__R2_INV_1 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y69__R3_BUF_0 (.A(tie_lo_T4Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y6__R0_BUF_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R0_INV_0 (.A(tie_lo_T4Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y6__R1_BUF_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R1_INV_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R2_INV_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y6__R2_INV_1 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y6__R3_BUF_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y70__R0_BUF_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R0_INV_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y70__R1_BUF_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R1_INV_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R2_INV_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y70__R2_INV_1 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y70__R3_BUF_0 (.A(tie_lo_T4Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y71__R0_BUF_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R0_INV_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y71__R1_BUF_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R1_INV_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R2_INV_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y71__R2_INV_1 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y71__R3_BUF_0 (.A(tie_lo_T4Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y72__R0_BUF_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R0_INV_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y72__R1_BUF_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R1_INV_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R2_INV_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y72__R2_INV_1 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y72__R3_BUF_0 (.A(tie_lo_T4Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y73__R0_BUF_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R0_INV_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y73__R1_BUF_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R1_INV_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R2_INV_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y73__R2_INV_1 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y73__R3_BUF_0 (.A(tie_lo_T4Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y74__R0_BUF_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R0_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y74__R1_BUF_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R1_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R2_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y74__R2_INV_1 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y74__R3_BUF_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y75__R0_BUF_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R0_INV_0 (.A(tie_lo_T4Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y75__R1_BUF_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R1_INV_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R2_INV_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y75__R2_INV_1 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y75__R3_BUF_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y76__R0_BUF_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R0_INV_0 (.A(tie_lo_T4Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y76__R1_BUF_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R1_INV_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R2_INV_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y76__R2_INV_1 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y76__R3_BUF_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y77__R0_BUF_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R0_INV_0 (.A(tie_lo_T4Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y77__R1_BUF_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R1_INV_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R2_INV_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y77__R2_INV_1 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y77__R3_BUF_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y78__R0_BUF_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R0_INV_0 (.A(tie_lo_T4Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y78__R1_BUF_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R1_INV_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R2_INV_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y78__R2_INV_1 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y78__R3_BUF_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y79__R0_BUF_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R0_INV_0 (.A(tie_lo_T4Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y79__R1_BUF_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R1_INV_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R2_INV_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y79__R2_INV_1 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y79__R3_BUF_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y7__R0_BUF_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R0_INV_0 (.A(tie_lo_T4Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y7__R1_BUF_0 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R1_INV_0 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R2_INV_0 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y7__R2_INV_1 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y7__R3_BUF_0 (.A(tie_lo_T4Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y80__R0_BUF_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R0_INV_0 (.A(tie_lo_T4Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y80__R1_BUF_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R1_INV_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R2_INV_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y80__R2_INV_1 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y80__R3_BUF_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y81__R0_BUF_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R0_INV_0 (.A(tie_lo_T4Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y81__R1_BUF_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R1_INV_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R2_INV_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y81__R2_INV_1 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y81__R3_BUF_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y82__R0_BUF_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R0_INV_0 (.A(tie_lo_T4Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y82__R1_BUF_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R1_INV_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R2_INV_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y82__R2_INV_1 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y82__R3_BUF_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y83__R0_BUF_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R0_INV_0 (.A(tie_lo_T4Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y83__R1_BUF_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R1_INV_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R2_INV_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y83__R2_INV_1 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y83__R3_BUF_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y84__R0_BUF_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R0_INV_0 (.A(tie_lo_T4Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y84__R1_BUF_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R1_INV_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R2_INV_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y84__R2_INV_1 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y84__R3_BUF_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y85__R0_BUF_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R0_INV_0 (.A(tie_lo_T4Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y85__R1_BUF_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R1_INV_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R2_INV_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y85__R2_INV_1 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y85__R3_BUF_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y86__R0_BUF_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R0_INV_0 (.A(tie_lo_T4Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y86__R1_BUF_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R1_INV_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R2_INV_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y86__R2_INV_1 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y86__R3_BUF_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y87__R0_BUF_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R0_INV_0 (.A(tie_lo_T4Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y87__R1_BUF_0 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R1_INV_0 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R2_INV_0 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y87__R2_INV_1 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y87__R3_BUF_0 (.A(tie_lo_T4Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y88__R0_BUF_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R0_INV_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y88__R1_BUF_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R1_INV_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R2_INV_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y88__R2_INV_1 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y88__R3_BUF_0 (.A(tie_lo_T4Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y89__R0_BUF_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R0_INV_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y89__R1_BUF_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R1_INV_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R2_INV_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y89__R2_INV_1 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y89__R3_BUF_0 (.A(tie_lo_T4Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y8__R0_BUF_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R0_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y8__R1_BUF_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R1_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R2_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y8__R2_INV_1 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y8__R3_BUF_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y9__R0_BUF_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R0_INV_0 (.A(tie_lo_T4Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y9__R1_BUF_0 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R1_INV_0 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T4Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R2_INV_0 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T4Y9__R2_INV_1 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T4Y9__R3_BUF_0 (.A(tie_lo_T4Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y0__R0_BUF_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R0_INV_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y0__R1_BUF_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R1_INV_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R2_INV_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y0__R2_INV_1 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y0__R3_BUF_0 (.A(tie_lo_T5Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y10__R0_BUF_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R0_INV_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y10__R1_BUF_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R1_INV_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R2_INV_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y10__R2_INV_1 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y10__R3_BUF_0 (.A(tie_lo_T5Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y11__R0_BUF_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R0_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y11__R1_BUF_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R1_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R2_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y11__R2_INV_1 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y11__R3_BUF_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y12__R0_BUF_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R0_INV_0 (.A(tie_lo_T5Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y12__R1_BUF_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R1_INV_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R2_INV_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y12__R2_INV_1 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y12__R3_BUF_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y13__R0_BUF_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R0_INV_0 (.A(tie_lo_T5Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y13__R1_BUF_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R1_INV_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R2_INV_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y13__R2_INV_1 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y13__R3_BUF_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y14__R0_BUF_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R0_INV_0 (.A(tie_lo_T5Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y14__R1_BUF_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R1_INV_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R2_INV_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y14__R2_INV_1 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y14__R3_BUF_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y15__R0_BUF_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R0_INV_0 (.A(tie_lo_T5Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y15__R1_BUF_0 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R1_INV_0 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R2_INV_0 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y15__R2_INV_1 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y15__R3_BUF_0 (.A(tie_lo_T5Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y16__R0_BUF_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R0_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y16__R1_BUF_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R1_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R2_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y16__R2_INV_1 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y16__R3_BUF_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y17__R0_BUF_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R0_INV_0 (.A(tie_lo_T5Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y17__R1_BUF_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R1_INV_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R2_INV_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y17__R2_INV_1 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y17__R3_BUF_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y18__R0_BUF_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R0_INV_0 (.A(tie_lo_T5Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y18__R1_BUF_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R1_INV_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R2_INV_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y18__R2_INV_1 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y18__R3_BUF_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y19__R0_BUF_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R0_INV_0 (.A(tie_lo_T5Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y19__R1_BUF_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R1_INV_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R2_INV_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y19__R2_INV_1 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y19__R3_BUF_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y1__R0_BUF_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R0_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y1__R1_BUF_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R1_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R2_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y1__R2_INV_1 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y1__R3_BUF_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y20__R0_BUF_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R0_INV_0 (.A(tie_lo_T5Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y20__R1_BUF_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R1_INV_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R2_INV_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y20__R2_INV_1 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y20__R3_BUF_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y21__R0_BUF_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R0_INV_0 (.A(tie_lo_T5Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y21__R1_BUF_0 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R1_INV_0 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R2_INV_0 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y21__R2_INV_1 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y21__R3_BUF_0 (.A(tie_lo_T5Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y22__R0_BUF_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R0_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y22__R1_BUF_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R1_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R2_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y22__R2_INV_1 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y22__R3_BUF_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y23__R0_BUF_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R0_INV_0 (.A(tie_lo_T5Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y23__R1_BUF_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R1_INV_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R2_INV_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y23__R2_INV_1 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y23__R3_BUF_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y24__R0_BUF_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R0_INV_0 (.A(tie_lo_T5Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y24__R1_BUF_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R1_INV_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R2_INV_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y24__R2_INV_1 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y24__R3_BUF_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y25__R0_BUF_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R0_INV_0 (.A(tie_lo_T5Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y25__R1_BUF_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R1_INV_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R2_INV_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y25__R2_INV_1 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y25__R3_BUF_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y26__R0_BUF_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R0_INV_0 (.A(tie_lo_T5Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y26__R1_BUF_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R1_INV_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R2_INV_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y26__R2_INV_1 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y26__R3_BUF_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y27__R0_BUF_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R0_INV_0 (.A(tie_lo_T5Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y27__R1_BUF_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R1_INV_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R2_INV_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y27__R2_INV_1 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y27__R3_BUF_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y28__R0_BUF_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R0_INV_0 (.A(tie_lo_T5Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y28__R1_BUF_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R1_INV_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R2_INV_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y28__R2_INV_1 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y28__R3_BUF_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y29__R0_BUF_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R0_INV_0 (.A(tie_lo_T5Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y29__R1_BUF_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R1_INV_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R2_INV_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y29__R2_INV_1 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y29__R3_BUF_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y2__R0_BUF_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R0_INV_0 (.A(tie_lo_T5Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y2__R1_BUF_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R1_INV_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R2_INV_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y2__R2_INV_1 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y2__R3_BUF_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y30__R0_BUF_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R0_INV_0 (.A(tie_lo_T5Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y30__R1_BUF_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R1_INV_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R2_INV_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y30__R2_INV_1 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y30__R3_BUF_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y31__R0_BUF_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R0_INV_0 (.A(tie_lo_T5Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y31__R1_BUF_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R1_INV_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R2_INV_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y31__R2_INV_1 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y31__R3_BUF_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y32__R0_BUF_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R0_INV_0 (.A(tie_lo_T5Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y32__R1_BUF_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R1_INV_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R2_INV_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y32__R2_INV_1 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y32__R3_BUF_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y33__R0_BUF_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R0_INV_0 (.A(tie_lo_T5Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y33__R1_BUF_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R1_INV_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R2_INV_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y33__R2_INV_1 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y33__R3_BUF_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y34__R0_BUF_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R0_INV_0 (.A(tie_lo_T5Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y34__R1_BUF_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R1_INV_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R2_INV_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y34__R2_INV_1 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y34__R3_BUF_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y35__R0_BUF_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R0_INV_0 (.A(tie_lo_T5Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y35__R1_BUF_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R1_INV_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R2_INV_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y35__R2_INV_1 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y35__R3_BUF_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y36__R0_BUF_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R0_INV_0 (.A(tie_lo_T5Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y36__R1_BUF_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R1_INV_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R2_INV_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y36__R2_INV_1 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y36__R3_BUF_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y37__R0_BUF_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R0_INV_0 (.A(tie_lo_T5Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y37__R1_BUF_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R1_INV_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R2_INV_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y37__R2_INV_1 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y37__R3_BUF_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y38__R0_BUF_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R0_INV_0 (.A(tie_lo_T5Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y38__R1_BUF_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R1_INV_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R2_INV_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y38__R2_INV_1 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y38__R3_BUF_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y39__R0_BUF_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R0_INV_0 (.A(tie_lo_T5Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y39__R1_BUF_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R1_INV_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R2_INV_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y39__R2_INV_1 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y39__R3_BUF_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y3__R0_BUF_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R0_INV_0 (.A(tie_lo_T5Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y3__R1_BUF_0 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R1_INV_0 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R2_INV_0 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y3__R2_INV_1 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y3__R3_BUF_0 (.A(tie_lo_T5Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y40__R0_BUF_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R0_INV_0 (.A(tie_lo_T5Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y40__R1_BUF_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R1_INV_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R2_INV_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y40__R2_INV_1 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y40__R3_BUF_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y41__R0_BUF_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R0_INV_0 (.A(tie_lo_T5Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y41__R1_BUF_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R1_INV_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R2_INV_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y41__R2_INV_1 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y41__R3_BUF_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y42__R0_BUF_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R0_INV_0 (.A(tie_lo_T5Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y42__R1_BUF_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R1_INV_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R2_INV_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y42__R2_INV_1 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y42__R3_BUF_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y43__R0_BUF_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R0_INV_0 (.A(tie_lo_T5Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y43__R1_BUF_0 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R1_INV_0 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R2_INV_0 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y43__R2_INV_1 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y43__R3_BUF_0 (.A(tie_lo_T5Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y44__R0_BUF_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R0_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y44__R1_BUF_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R1_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R2_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y44__R2_INV_1 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y44__R3_BUF_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y45__R0_BUF_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R0_INV_0 (.A(tie_lo_T5Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y45__R1_BUF_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R1_INV_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R2_INV_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y45__R2_INV_1 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y45__R3_BUF_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y46__R0_BUF_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R0_INV_0 (.A(tie_lo_T5Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y46__R1_BUF_0 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R1_INV_0 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R2_INV_0 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y46__R2_INV_1 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y46__R3_BUF_0 (.A(tie_lo_T5Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y47__R0_BUF_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R0_INV_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y47__R1_BUF_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R1_INV_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R2_INV_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y47__R2_INV_1 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y47__R3_BUF_0 (.A(tie_lo_T5Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y48__R0_BUF_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R0_INV_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y48__R1_BUF_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R1_INV_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R2_INV_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y48__R2_INV_1 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y48__R3_BUF_0 (.A(tie_lo_T5Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y49__R0_BUF_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R0_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y49__R1_BUF_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R1_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R2_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y49__R2_INV_1 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y49__R3_BUF_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y4__R0_BUF_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R0_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y4__R1_BUF_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R1_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R2_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y4__R2_INV_1 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y4__R3_BUF_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y50__R0_BUF_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R0_INV_0 (.A(tie_lo_T5Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y50__R1_BUF_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R1_INV_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R2_INV_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y50__R2_INV_1 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y50__R3_BUF_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y51__R0_BUF_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R0_INV_0 (.A(tie_lo_T5Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y51__R1_BUF_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R1_INV_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R2_INV_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y51__R2_INV_1 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y51__R3_BUF_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y52__R0_BUF_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R0_INV_0 (.A(tie_lo_T5Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y52__R1_BUF_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R1_INV_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R2_INV_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y52__R2_INV_1 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y52__R3_BUF_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y53__R0_BUF_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R0_INV_0 (.A(tie_lo_T5Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y53__R1_BUF_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R1_INV_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R2_INV_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y53__R2_INV_1 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y53__R3_BUF_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y54__R0_BUF_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R0_INV_0 (.A(tie_lo_T5Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y54__R1_BUF_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R1_INV_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R2_INV_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y54__R2_INV_1 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y54__R3_BUF_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y55__R0_BUF_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R0_INV_0 (.A(tie_lo_T5Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y55__R1_BUF_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R1_INV_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R2_INV_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y55__R2_INV_1 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y55__R3_BUF_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y56__R0_BUF_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R0_INV_0 (.A(tie_lo_T5Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y56__R1_BUF_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R1_INV_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R2_INV_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y56__R2_INV_1 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y56__R3_BUF_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y57__R0_BUF_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R0_INV_0 (.A(tie_lo_T5Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y57__R1_BUF_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R1_INV_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R2_INV_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y57__R2_INV_1 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y57__R3_BUF_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y58__R0_BUF_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R0_INV_0 (.A(tie_lo_T5Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y58__R1_BUF_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R1_INV_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R2_INV_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y58__R2_INV_1 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y58__R3_BUF_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y59__R0_BUF_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R0_INV_0 (.A(tie_lo_T5Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y59__R1_BUF_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R1_INV_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R2_INV_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y59__R2_INV_1 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y59__R3_BUF_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y5__R0_BUF_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R0_INV_0 (.A(tie_lo_T5Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y5__R1_BUF_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R1_INV_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R2_INV_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y5__R2_INV_1 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y5__R3_BUF_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y60__R0_BUF_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R0_INV_0 (.A(tie_lo_T5Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y60__R1_BUF_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R1_INV_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R2_INV_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y60__R2_INV_1 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y60__R3_BUF_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y61__R0_BUF_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R0_INV_0 (.A(tie_lo_T5Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y61__R1_BUF_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R1_INV_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R2_INV_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y61__R2_INV_1 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y61__R3_BUF_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y62__R0_BUF_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R0_INV_0 (.A(tie_lo_T5Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y62__R1_BUF_0 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R1_INV_0 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R2_INV_0 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y62__R2_INV_1 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y62__R3_BUF_0 (.A(tie_lo_T5Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y63__R0_BUF_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R0_INV_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y63__R1_BUF_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R1_INV_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R2_INV_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y63__R2_INV_1 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y63__R3_BUF_0 (.A(tie_lo_T5Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y64__R0_BUF_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R0_INV_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y64__R1_BUF_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R1_INV_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R2_INV_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y64__R2_INV_1 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y64__R3_BUF_0 (.A(tie_lo_T5Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y65__R0_BUF_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R0_INV_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y65__R1_BUF_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R1_INV_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R2_INV_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y65__R2_INV_1 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y65__R3_BUF_0 (.A(tie_lo_T5Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y66__R0_BUF_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R0_INV_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y66__R1_BUF_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R1_INV_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R2_INV_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y66__R2_INV_1 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y66__R3_BUF_0 (.A(tie_lo_T5Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y67__R0_BUF_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R0_INV_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y67__R1_BUF_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R1_INV_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R2_INV_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y67__R2_INV_1 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y67__R3_BUF_0 (.A(tie_lo_T5Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y68__R0_BUF_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R0_INV_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y68__R1_BUF_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R1_INV_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R2_INV_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y68__R2_INV_1 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y68__R3_BUF_0 (.A(tie_lo_T5Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y69__R0_BUF_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R0_INV_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y69__R1_BUF_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R1_INV_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R2_INV_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y69__R2_INV_1 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y69__R3_BUF_0 (.A(tie_lo_T5Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y6__R0_BUF_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R0_INV_0 (.A(tie_lo_T5Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y6__R1_BUF_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R1_INV_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R2_INV_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y6__R2_INV_1 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y6__R3_BUF_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y70__R0_BUF_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R0_INV_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y70__R1_BUF_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R1_INV_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R2_INV_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y70__R2_INV_1 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y70__R3_BUF_0 (.A(tie_lo_T5Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y71__R0_BUF_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R0_INV_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y71__R1_BUF_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R1_INV_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R2_INV_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y71__R2_INV_1 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y71__R3_BUF_0 (.A(tie_lo_T5Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y72__R0_BUF_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R0_INV_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y72__R1_BUF_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R1_INV_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R2_INV_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y72__R2_INV_1 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y72__R3_BUF_0 (.A(tie_lo_T5Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y73__R0_BUF_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R0_INV_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y73__R1_BUF_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R1_INV_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R2_INV_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y73__R2_INV_1 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y73__R3_BUF_0 (.A(tie_lo_T5Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y74__R0_BUF_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R0_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y74__R1_BUF_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R1_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R2_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y74__R2_INV_1 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y74__R3_BUF_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y75__R0_BUF_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R0_INV_0 (.A(tie_lo_T5Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y75__R1_BUF_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R1_INV_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R2_INV_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y75__R2_INV_1 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y75__R3_BUF_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y76__R0_BUF_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R0_INV_0 (.A(tie_lo_T5Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y76__R1_BUF_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R1_INV_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R2_INV_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y76__R2_INV_1 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y76__R3_BUF_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y77__R0_BUF_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R0_INV_0 (.A(tie_lo_T5Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y77__R1_BUF_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R1_INV_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R2_INV_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y77__R2_INV_1 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y77__R3_BUF_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y78__R0_BUF_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R0_INV_0 (.A(tie_lo_T5Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y78__R1_BUF_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R1_INV_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R2_INV_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y78__R2_INV_1 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y78__R3_BUF_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y79__R0_BUF_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R0_INV_0 (.A(tie_lo_T5Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y79__R1_BUF_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R1_INV_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R2_INV_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y79__R2_INV_1 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y79__R3_BUF_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y7__R0_BUF_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R0_INV_0 (.A(tie_lo_T5Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y7__R1_BUF_0 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R1_INV_0 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R2_INV_0 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y7__R2_INV_1 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y7__R3_BUF_0 (.A(tie_lo_T5Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y80__R0_BUF_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R0_INV_0 (.A(tie_lo_T5Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y80__R1_BUF_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R1_INV_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R2_INV_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y80__R2_INV_1 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y80__R3_BUF_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y81__R0_BUF_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R0_INV_0 (.A(tie_lo_T5Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y81__R1_BUF_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R1_INV_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R2_INV_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y81__R2_INV_1 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y81__R3_BUF_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y82__R0_BUF_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R0_INV_0 (.A(tie_lo_T5Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y82__R1_BUF_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R1_INV_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R2_INV_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y82__R2_INV_1 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y82__R3_BUF_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y83__R0_BUF_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R0_INV_0 (.A(tie_lo_T5Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y83__R1_BUF_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R1_INV_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R2_INV_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y83__R2_INV_1 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y83__R3_BUF_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y84__R0_BUF_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R0_INV_0 (.A(tie_lo_T5Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y84__R1_BUF_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R1_INV_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R2_INV_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y84__R2_INV_1 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y84__R3_BUF_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y85__R0_BUF_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R0_INV_0 (.A(tie_lo_T5Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y85__R1_BUF_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R1_INV_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R2_INV_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y85__R2_INV_1 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y85__R3_BUF_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y86__R0_BUF_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R0_INV_0 (.A(tie_lo_T5Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y86__R1_BUF_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R1_INV_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R2_INV_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y86__R2_INV_1 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y86__R3_BUF_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y87__R0_BUF_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R0_INV_0 (.A(tie_lo_T5Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y87__R1_BUF_0 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R1_INV_0 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R2_INV_0 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y87__R2_INV_1 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y87__R3_BUF_0 (.A(tie_lo_T5Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y88__R0_BUF_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R0_INV_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y88__R1_BUF_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R1_INV_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R2_INV_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y88__R2_INV_1 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y88__R3_BUF_0 (.A(tie_lo_T5Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y89__R0_BUF_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R0_INV_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y89__R1_BUF_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R1_INV_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R2_INV_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y89__R2_INV_1 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y89__R3_BUF_0 (.A(tie_lo_T5Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y8__R0_BUF_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R0_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y8__R1_BUF_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R1_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R2_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y8__R2_INV_1 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y8__R3_BUF_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y9__R0_BUF_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R0_INV_0 (.A(tie_lo_T5Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y9__R1_BUF_0 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R1_INV_0 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T5Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R2_INV_0 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T5Y9__R2_INV_1 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T5Y9__R3_BUF_0 (.A(tie_lo_T5Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y0__R0_BUF_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R0_INV_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y0__R1_BUF_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R1_INV_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R2_INV_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y0__R2_INV_1 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y0__R3_BUF_0 (.A(tie_lo_T6Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y10__R0_BUF_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R0_INV_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y10__R1_BUF_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R1_INV_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R2_INV_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y10__R2_INV_1 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y10__R3_BUF_0 (.A(tie_lo_T6Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y11__R0_BUF_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R0_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y11__R1_BUF_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R1_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R2_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y11__R2_INV_1 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y11__R3_BUF_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y12__R0_BUF_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R0_INV_0 (.A(tie_lo_T6Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y12__R1_BUF_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R1_INV_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R2_INV_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y12__R2_INV_1 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y12__R3_BUF_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y13__R0_BUF_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R0_INV_0 (.A(tie_lo_T6Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y13__R1_BUF_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R1_INV_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R2_INV_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y13__R2_INV_1 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y13__R3_BUF_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y14__R0_BUF_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R0_INV_0 (.A(tie_lo_T6Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y14__R1_BUF_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R1_INV_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R2_INV_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y14__R2_INV_1 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y14__R3_BUF_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y15__R0_BUF_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R0_INV_0 (.A(tie_lo_T6Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y15__R1_BUF_0 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R1_INV_0 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R2_INV_0 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y15__R2_INV_1 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y15__R3_BUF_0 (.A(tie_lo_T6Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y16__R0_BUF_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R0_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y16__R1_BUF_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R1_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R2_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y16__R2_INV_1 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y16__R3_BUF_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y17__R0_BUF_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R0_INV_0 (.A(tie_lo_T6Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y17__R1_BUF_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R1_INV_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R2_INV_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y17__R2_INV_1 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y17__R3_BUF_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y18__R0_BUF_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R0_INV_0 (.A(tie_lo_T6Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y18__R1_BUF_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R1_INV_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R2_INV_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y18__R2_INV_1 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y18__R3_BUF_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y19__R0_BUF_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R0_INV_0 (.A(tie_lo_T6Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y19__R1_BUF_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R1_INV_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R2_INV_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y19__R2_INV_1 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y19__R3_BUF_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y1__R0_BUF_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R0_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y1__R1_BUF_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R1_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R2_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y1__R2_INV_1 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y1__R3_BUF_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y20__R0_BUF_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R0_INV_0 (.A(tie_lo_T6Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y20__R1_BUF_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R1_INV_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R2_INV_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y20__R2_INV_1 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y20__R3_BUF_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y21__R0_BUF_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R0_INV_0 (.A(tie_lo_T6Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y21__R1_BUF_0 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R1_INV_0 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R2_INV_0 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y21__R2_INV_1 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y21__R3_BUF_0 (.A(tie_lo_T6Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y22__R0_BUF_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R0_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y22__R1_BUF_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R1_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R2_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y22__R2_INV_1 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y22__R3_BUF_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y23__R0_BUF_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R0_INV_0 (.A(tie_lo_T6Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y23__R1_BUF_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R1_INV_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R2_INV_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y23__R2_INV_1 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y23__R3_BUF_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y24__R0_BUF_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R0_INV_0 (.A(tie_lo_T6Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y24__R1_BUF_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R1_INV_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R2_INV_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y24__R2_INV_1 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y24__R3_BUF_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y25__R0_BUF_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R0_INV_0 (.A(tie_lo_T6Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y25__R1_BUF_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R1_INV_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R2_INV_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y25__R2_INV_1 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y25__R3_BUF_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y26__R0_BUF_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R0_INV_0 (.A(tie_lo_T6Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y26__R1_BUF_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R1_INV_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R2_INV_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y26__R2_INV_1 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y26__R3_BUF_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y27__R0_BUF_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R0_INV_0 (.A(tie_lo_T6Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y27__R1_BUF_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R1_INV_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R2_INV_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y27__R2_INV_1 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y27__R3_BUF_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y28__R0_BUF_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R0_INV_0 (.A(tie_lo_T6Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y28__R1_BUF_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R1_INV_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R2_INV_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y28__R2_INV_1 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y28__R3_BUF_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y29__R0_BUF_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R0_INV_0 (.A(tie_lo_T6Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y29__R1_BUF_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R1_INV_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R2_INV_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y29__R2_INV_1 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y29__R3_BUF_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y2__R0_BUF_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R0_INV_0 (.A(tie_lo_T6Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y2__R1_BUF_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R1_INV_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R2_INV_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y2__R2_INV_1 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y2__R3_BUF_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y30__R0_BUF_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R0_INV_0 (.A(tie_lo_T6Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y30__R1_BUF_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R1_INV_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R2_INV_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y30__R2_INV_1 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y30__R3_BUF_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y31__R0_BUF_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R0_INV_0 (.A(tie_lo_T6Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y31__R1_BUF_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R1_INV_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R2_INV_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y31__R2_INV_1 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y31__R3_BUF_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y32__R0_BUF_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R0_INV_0 (.A(tie_lo_T6Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y32__R1_BUF_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R1_INV_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R2_INV_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y32__R2_INV_1 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y32__R3_BUF_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y33__R0_BUF_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R0_INV_0 (.A(tie_lo_T6Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y33__R1_BUF_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R1_INV_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R2_INV_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y33__R2_INV_1 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y33__R3_BUF_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y34__R0_BUF_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R0_INV_0 (.A(tie_lo_T6Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y34__R1_BUF_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R1_INV_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R2_INV_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y34__R2_INV_1 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y34__R3_BUF_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y35__R0_BUF_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R0_INV_0 (.A(tie_lo_T6Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y35__R1_BUF_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R1_INV_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R2_INV_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y35__R2_INV_1 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y35__R3_BUF_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y36__R0_BUF_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R0_INV_0 (.A(tie_lo_T6Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y36__R1_BUF_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R1_INV_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R2_INV_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y36__R2_INV_1 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y36__R3_BUF_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y37__R0_BUF_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R0_INV_0 (.A(tie_lo_T6Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y37__R1_BUF_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R1_INV_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R2_INV_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y37__R2_INV_1 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y37__R3_BUF_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y38__R0_BUF_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R0_INV_0 (.A(tie_lo_T6Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y38__R1_BUF_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R1_INV_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R2_INV_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y38__R2_INV_1 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y38__R3_BUF_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y39__R0_BUF_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R0_INV_0 (.A(tie_lo_T6Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y39__R1_BUF_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R1_INV_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R2_INV_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y39__R2_INV_1 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y39__R3_BUF_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y3__R0_BUF_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R0_INV_0 (.A(tie_lo_T6Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y3__R1_BUF_0 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R1_INV_0 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R2_INV_0 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y3__R2_INV_1 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y3__R3_BUF_0 (.A(tie_lo_T6Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y40__R0_BUF_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R0_INV_0 (.A(tie_lo_T6Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y40__R1_BUF_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R1_INV_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R2_INV_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y40__R2_INV_1 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y40__R3_BUF_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y41__R0_BUF_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R0_INV_0 (.A(tie_lo_T6Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y41__R1_BUF_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R1_INV_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R2_INV_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y41__R2_INV_1 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y41__R3_BUF_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y42__R0_BUF_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R0_INV_0 (.A(tie_lo_T6Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y42__R1_BUF_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R1_INV_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R2_INV_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y42__R2_INV_1 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y42__R3_BUF_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y43__R0_BUF_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R0_INV_0 (.A(tie_lo_T6Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y43__R1_BUF_0 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R1_INV_0 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R2_INV_0 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y43__R2_INV_1 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y43__R3_BUF_0 (.A(tie_lo_T6Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y44__R0_BUF_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R0_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y44__R1_BUF_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R1_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R2_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y44__R2_INV_1 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y44__R3_BUF_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y45__R0_BUF_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R0_INV_0 (.A(tie_lo_T6Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y45__R1_BUF_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R1_INV_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R2_INV_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y45__R2_INV_1 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y45__R3_BUF_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y46__R0_BUF_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R0_INV_0 (.A(tie_lo_T6Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y46__R1_BUF_0 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R1_INV_0 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R2_INV_0 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y46__R2_INV_1 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y46__R3_BUF_0 (.A(tie_lo_T6Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y47__R0_BUF_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R0_INV_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y47__R1_BUF_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R1_INV_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R2_INV_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y47__R2_INV_1 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y47__R3_BUF_0 (.A(tie_lo_T6Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y48__R0_BUF_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R0_INV_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y48__R1_BUF_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R1_INV_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R2_INV_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y48__R2_INV_1 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y48__R3_BUF_0 (.A(tie_lo_T6Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y49__R0_BUF_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R0_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y49__R1_BUF_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R1_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R2_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y49__R2_INV_1 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y49__R3_BUF_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y4__R0_BUF_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R0_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y4__R1_BUF_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R1_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R2_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y4__R2_INV_1 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y4__R3_BUF_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y50__R0_BUF_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R0_INV_0 (.A(tie_lo_T6Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y50__R1_BUF_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R1_INV_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R2_INV_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y50__R2_INV_1 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y50__R3_BUF_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y51__R0_BUF_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R0_INV_0 (.A(tie_lo_T6Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y51__R1_BUF_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R1_INV_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R2_INV_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y51__R2_INV_1 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y51__R3_BUF_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y52__R0_BUF_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R0_INV_0 (.A(tie_lo_T6Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y52__R1_BUF_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R1_INV_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R2_INV_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y52__R2_INV_1 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y52__R3_BUF_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y53__R0_BUF_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R0_INV_0 (.A(tie_lo_T6Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y53__R1_BUF_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R1_INV_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R2_INV_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y53__R2_INV_1 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y53__R3_BUF_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y54__R0_BUF_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R0_INV_0 (.A(tie_lo_T6Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y54__R1_BUF_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R1_INV_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R2_INV_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y54__R2_INV_1 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y54__R3_BUF_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y55__R0_BUF_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R0_INV_0 (.A(tie_lo_T6Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y55__R1_BUF_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R1_INV_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R2_INV_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y55__R2_INV_1 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y55__R3_BUF_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y56__R0_BUF_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R0_INV_0 (.A(tie_lo_T6Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y56__R1_BUF_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R1_INV_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R2_INV_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y56__R2_INV_1 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y56__R3_BUF_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y57__R0_BUF_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R0_INV_0 (.A(tie_lo_T6Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y57__R1_BUF_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R1_INV_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R2_INV_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y57__R2_INV_1 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y57__R3_BUF_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y58__R0_BUF_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R0_INV_0 (.A(tie_lo_T6Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y58__R1_BUF_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R1_INV_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R2_INV_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y58__R2_INV_1 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y58__R3_BUF_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y59__R0_BUF_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R0_INV_0 (.A(tie_lo_T6Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y59__R1_BUF_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R1_INV_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R2_INV_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y59__R2_INV_1 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y59__R3_BUF_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y5__R0_BUF_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R0_INV_0 (.A(tie_lo_T6Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y5__R1_BUF_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R1_INV_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R2_INV_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y5__R2_INV_1 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y5__R3_BUF_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y60__R0_BUF_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R0_INV_0 (.A(tie_lo_T6Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y60__R1_BUF_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R1_INV_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R2_INV_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y60__R2_INV_1 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y60__R3_BUF_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y61__R0_BUF_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R0_INV_0 (.A(tie_lo_T6Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y61__R1_BUF_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R1_INV_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R2_INV_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y61__R2_INV_1 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y61__R3_BUF_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y62__R0_BUF_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R0_INV_0 (.A(tie_lo_T6Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y62__R1_BUF_0 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R1_INV_0 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R2_INV_0 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y62__R2_INV_1 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y62__R3_BUF_0 (.A(tie_lo_T6Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y63__R0_BUF_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R0_INV_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y63__R1_BUF_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R1_INV_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R2_INV_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y63__R2_INV_1 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y63__R3_BUF_0 (.A(tie_lo_T6Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y64__R0_BUF_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R0_INV_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y64__R1_BUF_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R1_INV_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R2_INV_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y64__R2_INV_1 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y64__R3_BUF_0 (.A(tie_lo_T6Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y65__R0_BUF_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R0_INV_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y65__R1_BUF_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R1_INV_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R2_INV_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y65__R2_INV_1 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y65__R3_BUF_0 (.A(tie_lo_T6Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y66__R0_BUF_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R0_INV_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y66__R1_BUF_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R1_INV_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R2_INV_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y66__R2_INV_1 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y66__R3_BUF_0 (.A(tie_lo_T6Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y67__R0_BUF_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R0_INV_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y67__R1_BUF_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R1_INV_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R2_INV_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y67__R2_INV_1 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y67__R3_BUF_0 (.A(tie_lo_T6Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y68__R0_BUF_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R0_INV_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y68__R1_BUF_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R1_INV_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R2_INV_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y68__R2_INV_1 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y68__R3_BUF_0 (.A(tie_lo_T6Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y69__R0_BUF_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R0_INV_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y69__R1_BUF_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R1_INV_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R2_INV_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y69__R2_INV_1 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y69__R3_BUF_0 (.A(tie_lo_T6Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y6__R0_BUF_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R0_INV_0 (.A(tie_lo_T6Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y6__R1_BUF_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R1_INV_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R2_INV_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y6__R2_INV_1 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y6__R3_BUF_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y70__R0_BUF_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R0_INV_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y70__R1_BUF_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R1_INV_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R2_INV_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y70__R2_INV_1 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y70__R3_BUF_0 (.A(tie_lo_T6Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y71__R0_BUF_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R0_INV_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y71__R1_BUF_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R1_INV_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R2_INV_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y71__R2_INV_1 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y71__R3_BUF_0 (.A(tie_lo_T6Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y72__R0_BUF_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R0_INV_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y72__R1_BUF_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R1_INV_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R2_INV_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y72__R2_INV_1 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y72__R3_BUF_0 (.A(tie_lo_T6Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y73__R0_BUF_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R0_INV_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y73__R1_BUF_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R1_INV_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R2_INV_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y73__R2_INV_1 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y73__R3_BUF_0 (.A(tie_lo_T6Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y74__R0_BUF_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R0_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y74__R1_BUF_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R1_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R2_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y74__R2_INV_1 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y74__R3_BUF_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y75__R0_BUF_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R0_INV_0 (.A(tie_lo_T6Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y75__R1_BUF_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R1_INV_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R2_INV_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y75__R2_INV_1 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y75__R3_BUF_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y76__R0_BUF_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R0_INV_0 (.A(tie_lo_T6Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y76__R1_BUF_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R1_INV_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R2_INV_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y76__R2_INV_1 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y76__R3_BUF_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y77__R0_BUF_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R0_INV_0 (.A(tie_lo_T6Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y77__R1_BUF_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R1_INV_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R2_INV_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y77__R2_INV_1 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y77__R3_BUF_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y78__R0_BUF_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R0_INV_0 (.A(tie_lo_T6Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y78__R1_BUF_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R1_INV_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R2_INV_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y78__R2_INV_1 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y78__R3_BUF_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y79__R0_BUF_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R0_INV_0 (.A(tie_lo_T6Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y79__R1_BUF_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R1_INV_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R2_INV_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y79__R2_INV_1 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y79__R3_BUF_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y7__R0_BUF_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R0_INV_0 (.A(tie_lo_T6Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y7__R1_BUF_0 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R1_INV_0 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R2_INV_0 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y7__R2_INV_1 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y7__R3_BUF_0 (.A(tie_lo_T6Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y80__R0_BUF_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R0_INV_0 (.A(tie_lo_T6Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y80__R1_BUF_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R1_INV_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R2_INV_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y80__R2_INV_1 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y80__R3_BUF_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y81__R0_BUF_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R0_INV_0 (.A(tie_lo_T6Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y81__R1_BUF_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R1_INV_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R2_INV_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y81__R2_INV_1 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y81__R3_BUF_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y82__R0_BUF_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R0_INV_0 (.A(tie_lo_T6Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y82__R1_BUF_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R1_INV_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R2_INV_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y82__R2_INV_1 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y82__R3_BUF_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y83__R0_BUF_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R0_INV_0 (.A(tie_lo_T6Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y83__R1_BUF_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R1_INV_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R2_INV_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y83__R2_INV_1 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y83__R3_BUF_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y84__R0_BUF_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R0_INV_0 (.A(tie_lo_T6Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y84__R1_BUF_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R1_INV_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R2_INV_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y84__R2_INV_1 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y84__R3_BUF_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y85__R0_BUF_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R0_INV_0 (.A(tie_lo_T6Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y85__R1_BUF_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R1_INV_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R2_INV_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y85__R2_INV_1 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y85__R3_BUF_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y86__R0_BUF_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R0_INV_0 (.A(tie_lo_T6Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y86__R1_BUF_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R1_INV_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R2_INV_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y86__R2_INV_1 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y86__R3_BUF_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y87__R0_BUF_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R0_INV_0 (.A(tie_lo_T6Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y87__R1_BUF_0 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R1_INV_0 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R2_INV_0 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y87__R2_INV_1 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y87__R3_BUF_0 (.A(tie_lo_T6Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y88__R0_BUF_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R0_INV_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y88__R1_BUF_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R1_INV_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R2_INV_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y88__R2_INV_1 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y88__R3_BUF_0 (.A(tie_lo_T6Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y89__R0_BUF_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R0_INV_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y89__R1_BUF_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R1_INV_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R2_INV_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y89__R2_INV_1 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y89__R3_BUF_0 (.A(tie_lo_T6Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y8__R0_BUF_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R0_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y8__R1_BUF_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R1_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R2_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y8__R2_INV_1 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y8__R3_BUF_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y9__R0_BUF_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R0_INV_0 (.A(tie_lo_T6Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y9__R1_BUF_0 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R1_INV_0 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T6Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R2_INV_0 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T6Y9__R2_INV_1 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T6Y9__R3_BUF_0 (.A(tie_lo_T6Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y0__R0_BUF_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R0_INV_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y0__R1_BUF_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R1_INV_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R2_INV_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y0__R2_INV_1 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y0__R3_BUF_0 (.A(tie_lo_T7Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y10__R0_BUF_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R0_INV_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y10__R1_BUF_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R1_INV_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R2_INV_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y10__R2_INV_1 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y10__R3_BUF_0 (.A(tie_lo_T7Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y11__R0_BUF_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R0_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y11__R1_BUF_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R1_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R2_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y11__R2_INV_1 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y11__R3_BUF_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y12__R0_BUF_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R0_INV_0 (.A(tie_lo_T7Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y12__R1_BUF_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R1_INV_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R2_INV_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y12__R2_INV_1 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y12__R3_BUF_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y13__R0_BUF_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R0_INV_0 (.A(tie_lo_T7Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y13__R1_BUF_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R1_INV_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R2_INV_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y13__R2_INV_1 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y13__R3_BUF_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y14__R0_BUF_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R0_INV_0 (.A(tie_lo_T7Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y14__R1_BUF_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R1_INV_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R2_INV_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y14__R2_INV_1 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y14__R3_BUF_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y15__R0_BUF_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R0_INV_0 (.A(tie_lo_T7Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y15__R1_BUF_0 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R1_INV_0 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R2_INV_0 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y15__R2_INV_1 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y15__R3_BUF_0 (.A(tie_lo_T7Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y16__R0_BUF_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R0_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y16__R1_BUF_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R1_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R2_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y16__R2_INV_1 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y16__R3_BUF_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y17__R0_BUF_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R0_INV_0 (.A(tie_lo_T7Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y17__R1_BUF_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R1_INV_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R2_INV_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y17__R2_INV_1 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y17__R3_BUF_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y18__R0_BUF_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R0_INV_0 (.A(tie_lo_T7Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y18__R1_BUF_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R1_INV_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R2_INV_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y18__R2_INV_1 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y18__R3_BUF_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y19__R0_BUF_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R0_INV_0 (.A(tie_lo_T7Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y19__R1_BUF_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R1_INV_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R2_INV_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y19__R2_INV_1 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y19__R3_BUF_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y1__R0_BUF_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R0_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y1__R1_BUF_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R1_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R2_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y1__R2_INV_1 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y1__R3_BUF_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y20__R0_BUF_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R0_INV_0 (.A(tie_lo_T7Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y20__R1_BUF_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R1_INV_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R2_INV_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y20__R2_INV_1 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y20__R3_BUF_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y21__R0_BUF_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R0_INV_0 (.A(tie_lo_T7Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y21__R1_BUF_0 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R1_INV_0 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R2_INV_0 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y21__R2_INV_1 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y21__R3_BUF_0 (.A(tie_lo_T7Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y22__R0_BUF_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R0_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y22__R1_BUF_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R1_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R2_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y22__R2_INV_1 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y22__R3_BUF_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y23__R0_BUF_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R0_INV_0 (.A(tie_lo_T7Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y23__R1_BUF_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R1_INV_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R2_INV_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y23__R2_INV_1 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y23__R3_BUF_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y24__R0_BUF_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R0_INV_0 (.A(tie_lo_T7Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y24__R1_BUF_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R1_INV_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R2_INV_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y24__R2_INV_1 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y24__R3_BUF_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y25__R0_BUF_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R0_INV_0 (.A(tie_lo_T7Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y25__R1_BUF_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R1_INV_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R2_INV_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y25__R2_INV_1 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y25__R3_BUF_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y26__R0_BUF_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R0_INV_0 (.A(tie_lo_T7Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y26__R1_BUF_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R1_INV_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R2_INV_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y26__R2_INV_1 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y26__R3_BUF_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y27__R0_BUF_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R0_INV_0 (.A(tie_lo_T7Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y27__R1_BUF_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R1_INV_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R2_INV_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y27__R2_INV_1 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y27__R3_BUF_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y28__R0_BUF_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R0_INV_0 (.A(tie_lo_T7Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y28__R1_BUF_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R1_INV_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R2_INV_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y28__R2_INV_1 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y28__R3_BUF_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y29__R0_BUF_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R0_INV_0 (.A(tie_lo_T7Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y29__R1_BUF_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R1_INV_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R2_INV_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y29__R2_INV_1 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y29__R3_BUF_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y2__R0_BUF_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R0_INV_0 (.A(tie_lo_T7Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y2__R1_BUF_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R1_INV_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R2_INV_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y2__R2_INV_1 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y2__R3_BUF_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y30__R0_BUF_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R0_INV_0 (.A(tie_lo_T7Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y30__R1_BUF_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R1_INV_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R2_INV_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y30__R2_INV_1 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y30__R3_BUF_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y31__R0_BUF_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R0_INV_0 (.A(tie_lo_T7Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y31__R1_BUF_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R1_INV_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R2_INV_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y31__R2_INV_1 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y31__R3_BUF_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y32__R0_BUF_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R0_INV_0 (.A(tie_lo_T7Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y32__R1_BUF_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R1_INV_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R2_INV_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y32__R2_INV_1 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y32__R3_BUF_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y33__R0_BUF_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R0_INV_0 (.A(tie_lo_T7Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y33__R1_BUF_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R1_INV_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R2_INV_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y33__R2_INV_1 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y33__R3_BUF_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y34__R0_BUF_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R0_INV_0 (.A(tie_lo_T7Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y34__R1_BUF_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R1_INV_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R2_INV_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y34__R2_INV_1 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y34__R3_BUF_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y35__R0_BUF_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R0_INV_0 (.A(tie_lo_T7Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y35__R1_BUF_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R1_INV_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R2_INV_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y35__R2_INV_1 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y35__R3_BUF_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y36__R0_BUF_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R0_INV_0 (.A(tie_lo_T7Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y36__R1_BUF_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R1_INV_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R2_INV_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y36__R2_INV_1 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y36__R3_BUF_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y37__R0_BUF_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R0_INV_0 (.A(tie_lo_T7Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y37__R1_BUF_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R1_INV_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R2_INV_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y37__R2_INV_1 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y37__R3_BUF_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y38__R0_BUF_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R0_INV_0 (.A(tie_lo_T7Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y38__R1_BUF_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R1_INV_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R2_INV_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y38__R2_INV_1 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y38__R3_BUF_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y39__R0_BUF_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R0_INV_0 (.A(tie_lo_T7Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y39__R1_BUF_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R1_INV_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R2_INV_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y39__R2_INV_1 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y39__R3_BUF_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y3__R0_BUF_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R0_INV_0 (.A(tie_lo_T7Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y3__R1_BUF_0 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R1_INV_0 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R2_INV_0 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y3__R2_INV_1 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y3__R3_BUF_0 (.A(tie_lo_T7Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y40__R0_BUF_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R0_INV_0 (.A(tie_lo_T7Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y40__R1_BUF_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R1_INV_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R2_INV_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y40__R2_INV_1 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y40__R3_BUF_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y41__R0_BUF_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R0_INV_0 (.A(tie_lo_T7Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y41__R1_BUF_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R1_INV_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R2_INV_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y41__R2_INV_1 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y41__R3_BUF_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y42__R0_BUF_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R0_INV_0 (.A(tie_lo_T7Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y42__R1_BUF_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R1_INV_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R2_INV_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y42__R2_INV_1 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y42__R3_BUF_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y43__R0_BUF_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R0_INV_0 (.A(tie_lo_T7Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y43__R1_BUF_0 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R1_INV_0 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R2_INV_0 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y43__R2_INV_1 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y43__R3_BUF_0 (.A(tie_lo_T7Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y44__R0_BUF_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R0_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y44__R1_BUF_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R1_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R2_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y44__R2_INV_1 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y44__R3_BUF_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y45__R0_BUF_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R0_INV_0 (.A(tie_lo_T7Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y45__R1_BUF_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R1_INV_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R2_INV_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y45__R2_INV_1 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y45__R3_BUF_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y46__R0_BUF_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R0_INV_0 (.A(tie_lo_T7Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y46__R1_BUF_0 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R1_INV_0 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R2_INV_0 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y46__R2_INV_1 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y46__R3_BUF_0 (.A(tie_lo_T7Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y47__R0_BUF_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R0_INV_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y47__R1_BUF_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R1_INV_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R2_INV_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y47__R2_INV_1 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y47__R3_BUF_0 (.A(tie_lo_T7Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y48__R0_BUF_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R0_INV_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y48__R1_BUF_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R1_INV_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R2_INV_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y48__R2_INV_1 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y48__R3_BUF_0 (.A(tie_lo_T7Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y49__R0_BUF_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R0_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y49__R1_BUF_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R1_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R2_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y49__R2_INV_1 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y49__R3_BUF_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y4__R0_BUF_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R0_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y4__R1_BUF_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R1_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R2_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y4__R2_INV_1 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y4__R3_BUF_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y50__R0_BUF_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R0_INV_0 (.A(tie_lo_T7Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y50__R1_BUF_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R1_INV_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R2_INV_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y50__R2_INV_1 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y50__R3_BUF_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y51__R0_BUF_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R0_INV_0 (.A(tie_lo_T7Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y51__R1_BUF_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R1_INV_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R2_INV_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y51__R2_INV_1 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y51__R3_BUF_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y52__R0_BUF_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R0_INV_0 (.A(tie_lo_T7Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y52__R1_BUF_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R1_INV_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R2_INV_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y52__R2_INV_1 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y52__R3_BUF_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y53__R0_BUF_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R0_INV_0 (.A(tie_lo_T7Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y53__R1_BUF_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R1_INV_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R2_INV_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y53__R2_INV_1 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y53__R3_BUF_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y54__R0_BUF_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R0_INV_0 (.A(tie_lo_T7Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y54__R1_BUF_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R1_INV_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R2_INV_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y54__R2_INV_1 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y54__R3_BUF_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y55__R0_BUF_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R0_INV_0 (.A(tie_lo_T7Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y55__R1_BUF_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R1_INV_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R2_INV_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y55__R2_INV_1 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y55__R3_BUF_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y56__R0_BUF_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R0_INV_0 (.A(tie_lo_T7Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y56__R1_BUF_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R1_INV_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R2_INV_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y56__R2_INV_1 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y56__R3_BUF_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y57__R0_BUF_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R0_INV_0 (.A(tie_lo_T7Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y57__R1_BUF_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R1_INV_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R2_INV_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y57__R2_INV_1 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y57__R3_BUF_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y58__R0_BUF_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R0_INV_0 (.A(tie_lo_T7Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y58__R1_BUF_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R1_INV_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R2_INV_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y58__R2_INV_1 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y58__R3_BUF_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y59__R0_BUF_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R0_INV_0 (.A(tie_lo_T7Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y59__R1_BUF_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R1_INV_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R2_INV_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y59__R2_INV_1 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y59__R3_BUF_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y5__R0_BUF_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R0_INV_0 (.A(tie_lo_T7Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y5__R1_BUF_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R1_INV_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R2_INV_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y5__R2_INV_1 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y5__R3_BUF_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y60__R0_BUF_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R0_INV_0 (.A(tie_lo_T7Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y60__R1_BUF_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R1_INV_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R2_INV_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y60__R2_INV_1 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y60__R3_BUF_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y61__R0_BUF_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R0_INV_0 (.A(tie_lo_T7Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y61__R1_BUF_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R1_INV_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R2_INV_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y61__R2_INV_1 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y61__R3_BUF_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y62__R0_BUF_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R0_INV_0 (.A(tie_lo_T7Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y62__R1_BUF_0 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R1_INV_0 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R2_INV_0 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y62__R2_INV_1 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y62__R3_BUF_0 (.A(tie_lo_T7Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y63__R0_BUF_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R0_INV_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y63__R1_BUF_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R1_INV_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R2_INV_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y63__R2_INV_1 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y63__R3_BUF_0 (.A(tie_lo_T7Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y64__R0_BUF_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R0_INV_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y64__R1_BUF_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R1_INV_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R2_INV_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y64__R2_INV_1 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y64__R3_BUF_0 (.A(tie_lo_T7Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y65__R0_BUF_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R0_INV_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y65__R1_BUF_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R1_INV_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R2_INV_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y65__R2_INV_1 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y65__R3_BUF_0 (.A(tie_lo_T7Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y66__R0_BUF_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R0_INV_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y66__R1_BUF_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R1_INV_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R2_INV_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y66__R2_INV_1 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y66__R3_BUF_0 (.A(tie_lo_T7Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y67__R0_BUF_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R0_INV_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y67__R1_BUF_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R1_INV_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R2_INV_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y67__R2_INV_1 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y67__R3_BUF_0 (.A(tie_lo_T7Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y68__R0_BUF_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R0_INV_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y68__R1_BUF_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R1_INV_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R2_INV_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y68__R2_INV_1 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y68__R3_BUF_0 (.A(tie_lo_T7Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y69__R0_BUF_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R0_INV_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y69__R1_BUF_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R1_INV_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R2_INV_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y69__R2_INV_1 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y69__R3_BUF_0 (.A(tie_lo_T7Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y6__R0_BUF_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R0_INV_0 (.A(tie_lo_T7Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y6__R1_BUF_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R1_INV_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R2_INV_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y6__R2_INV_1 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y6__R3_BUF_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y70__R0_BUF_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R0_INV_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y70__R1_BUF_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R1_INV_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R2_INV_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y70__R2_INV_1 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y70__R3_BUF_0 (.A(tie_lo_T7Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y71__R0_BUF_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R0_INV_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y71__R1_BUF_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R1_INV_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R2_INV_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y71__R2_INV_1 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y71__R3_BUF_0 (.A(tie_lo_T7Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y72__R0_BUF_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R0_INV_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y72__R1_BUF_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R1_INV_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R2_INV_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y72__R2_INV_1 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y72__R3_BUF_0 (.A(tie_lo_T7Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y73__R0_BUF_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R0_INV_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y73__R1_BUF_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R1_INV_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R2_INV_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y73__R2_INV_1 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y73__R3_BUF_0 (.A(tie_lo_T7Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y74__R0_BUF_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R0_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y74__R1_BUF_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R1_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R2_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y74__R2_INV_1 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y74__R3_BUF_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y75__R0_BUF_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R0_INV_0 (.A(tie_lo_T7Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y75__R1_BUF_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R1_INV_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R2_INV_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y75__R2_INV_1 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y75__R3_BUF_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y76__R0_BUF_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R0_INV_0 (.A(tie_lo_T7Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y76__R1_BUF_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R1_INV_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R2_INV_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y76__R2_INV_1 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y76__R3_BUF_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y77__R0_BUF_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R0_INV_0 (.A(tie_lo_T7Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y77__R1_BUF_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R1_INV_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R2_INV_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y77__R2_INV_1 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y77__R3_BUF_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y78__R0_BUF_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R0_INV_0 (.A(tie_lo_T7Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y78__R1_BUF_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R1_INV_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R2_INV_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y78__R2_INV_1 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y78__R3_BUF_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y79__R0_BUF_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R0_INV_0 (.A(tie_lo_T7Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y79__R1_BUF_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R1_INV_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R2_INV_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y79__R2_INV_1 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y79__R3_BUF_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y7__R0_BUF_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R0_INV_0 (.A(tie_lo_T7Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y7__R1_BUF_0 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R1_INV_0 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R2_INV_0 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y7__R2_INV_1 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y7__R3_BUF_0 (.A(tie_lo_T7Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y80__R0_BUF_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R0_INV_0 (.A(tie_lo_T7Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y80__R1_BUF_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R1_INV_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R2_INV_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y80__R2_INV_1 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y80__R3_BUF_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y81__R0_BUF_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R0_INV_0 (.A(tie_lo_T7Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y81__R1_BUF_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R1_INV_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R2_INV_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y81__R2_INV_1 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y81__R3_BUF_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y82__R0_BUF_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R0_INV_0 (.A(tie_lo_T7Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y82__R1_BUF_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R1_INV_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R2_INV_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y82__R2_INV_1 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y82__R3_BUF_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y83__R0_BUF_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R0_INV_0 (.A(tie_lo_T7Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y83__R1_BUF_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R1_INV_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R2_INV_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y83__R2_INV_1 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y83__R3_BUF_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y84__R0_BUF_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R0_INV_0 (.A(tie_lo_T7Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y84__R1_BUF_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R1_INV_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R2_INV_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y84__R2_INV_1 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y84__R3_BUF_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y85__R0_BUF_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R0_INV_0 (.A(tie_lo_T7Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y85__R1_BUF_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R1_INV_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R2_INV_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y85__R2_INV_1 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y85__R3_BUF_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y86__R0_BUF_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R0_INV_0 (.A(tie_lo_T7Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y86__R1_BUF_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R1_INV_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R2_INV_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y86__R2_INV_1 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y86__R3_BUF_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y87__R0_BUF_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R0_INV_0 (.A(tie_lo_T7Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y87__R1_BUF_0 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R1_INV_0 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R2_INV_0 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y87__R2_INV_1 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y87__R3_BUF_0 (.A(tie_lo_T7Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y88__R0_BUF_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R0_INV_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y88__R1_BUF_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R1_INV_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R2_INV_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y88__R2_INV_1 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y88__R3_BUF_0 (.A(tie_lo_T7Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y89__R0_BUF_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R0_INV_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y89__R1_BUF_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R1_INV_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R2_INV_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y89__R2_INV_1 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y89__R3_BUF_0 (.A(tie_lo_T7Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y8__R0_BUF_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R0_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y8__R1_BUF_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R1_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R2_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y8__R2_INV_1 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y8__R3_BUF_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y9__R0_BUF_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R0_INV_0 (.A(tie_lo_T7Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y9__R1_BUF_0 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R1_INV_0 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T7Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R2_INV_0 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T7Y9__R2_INV_1 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T7Y9__R3_BUF_0 (.A(tie_lo_T7Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y0__R0_BUF_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R0_INV_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y0__R1_BUF_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R1_INV_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R2_INV_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y0__R2_INV_1 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y0__R3_BUF_0 (.A(tie_lo_T8Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y10__R0_BUF_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R0_INV_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y10__R1_BUF_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R1_INV_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R2_INV_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y10__R2_INV_1 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y10__R3_BUF_0 (.A(tie_lo_T8Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y11__R0_BUF_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R0_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y11__R1_BUF_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R1_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R2_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y11__R2_INV_1 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y11__R3_BUF_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y12__R0_BUF_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R0_INV_0 (.A(tie_lo_T8Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y12__R1_BUF_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R1_INV_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R2_INV_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y12__R2_INV_1 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y12__R3_BUF_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y13__R0_BUF_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R0_INV_0 (.A(tie_lo_T8Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y13__R1_BUF_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R1_INV_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R2_INV_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y13__R2_INV_1 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y13__R3_BUF_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y14__R0_BUF_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R0_INV_0 (.A(tie_lo_T8Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y14__R1_BUF_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R1_INV_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R2_INV_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y14__R2_INV_1 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y14__R3_BUF_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y15__R0_BUF_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R0_INV_0 (.A(tie_lo_T8Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y15__R1_BUF_0 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R1_INV_0 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R2_INV_0 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y15__R2_INV_1 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y15__R3_BUF_0 (.A(tie_lo_T8Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y16__R0_BUF_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R0_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y16__R1_BUF_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R1_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R2_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y16__R2_INV_1 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y16__R3_BUF_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y17__R0_BUF_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R0_INV_0 (.A(tie_lo_T8Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y17__R1_BUF_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R1_INV_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R2_INV_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y17__R2_INV_1 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y17__R3_BUF_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y18__R0_BUF_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R0_INV_0 (.A(tie_lo_T8Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y18__R1_BUF_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R1_INV_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R2_INV_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y18__R2_INV_1 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y18__R3_BUF_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y19__R0_BUF_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R0_INV_0 (.A(tie_lo_T8Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y19__R1_BUF_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R1_INV_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R2_INV_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y19__R2_INV_1 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y19__R3_BUF_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y1__R0_BUF_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R0_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y1__R1_BUF_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R1_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R2_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y1__R2_INV_1 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y1__R3_BUF_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y20__R0_BUF_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R0_INV_0 (.A(tie_lo_T8Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y20__R1_BUF_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R1_INV_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R2_INV_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y20__R2_INV_1 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y20__R3_BUF_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y21__R0_BUF_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R0_INV_0 (.A(tie_lo_T8Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y21__R1_BUF_0 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R1_INV_0 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R2_INV_0 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y21__R2_INV_1 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y21__R3_BUF_0 (.A(tie_lo_T8Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y22__R0_BUF_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R0_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y22__R1_BUF_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R1_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R2_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y22__R2_INV_1 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y22__R3_BUF_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y23__R0_BUF_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R0_INV_0 (.A(tie_lo_T8Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y23__R1_BUF_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R1_INV_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R2_INV_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y23__R2_INV_1 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y23__R3_BUF_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y24__R0_BUF_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R0_INV_0 (.A(tie_lo_T8Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y24__R1_BUF_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R1_INV_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R2_INV_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y24__R2_INV_1 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y24__R3_BUF_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y25__R0_BUF_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R0_INV_0 (.A(tie_lo_T8Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y25__R1_BUF_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R1_INV_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R2_INV_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y25__R2_INV_1 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y25__R3_BUF_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y26__R0_BUF_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R0_INV_0 (.A(tie_lo_T8Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y26__R1_BUF_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R1_INV_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R2_INV_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y26__R2_INV_1 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y26__R3_BUF_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y27__R0_BUF_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R0_INV_0 (.A(tie_lo_T8Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y27__R1_BUF_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R1_INV_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R2_INV_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y27__R2_INV_1 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y27__R3_BUF_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y28__R0_BUF_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R0_INV_0 (.A(tie_lo_T8Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y28__R1_BUF_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R1_INV_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R2_INV_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y28__R2_INV_1 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y28__R3_BUF_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y29__R0_BUF_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R0_INV_0 (.A(tie_lo_T8Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y29__R1_BUF_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R1_INV_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R2_INV_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y29__R2_INV_1 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y29__R3_BUF_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y2__R0_BUF_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R0_INV_0 (.A(tie_lo_T8Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y2__R1_BUF_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R1_INV_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R2_INV_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y2__R2_INV_1 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y2__R3_BUF_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y30__R0_BUF_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R0_INV_0 (.A(tie_lo_T8Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y30__R1_BUF_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R1_INV_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R2_INV_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y30__R2_INV_1 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y30__R3_BUF_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y31__R0_BUF_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R0_INV_0 (.A(tie_lo_T8Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y31__R1_BUF_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R1_INV_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R2_INV_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y31__R2_INV_1 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y31__R3_BUF_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y32__R0_BUF_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R0_INV_0 (.A(tie_lo_T8Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y32__R1_BUF_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R1_INV_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R2_INV_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y32__R2_INV_1 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y32__R3_BUF_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y33__R0_BUF_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R0_INV_0 (.A(tie_lo_T8Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y33__R1_BUF_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R1_INV_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R2_INV_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y33__R2_INV_1 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y33__R3_BUF_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y34__R0_BUF_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R0_INV_0 (.A(tie_lo_T8Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y34__R1_BUF_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R1_INV_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R2_INV_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y34__R2_INV_1 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y34__R3_BUF_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y35__R0_BUF_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R0_INV_0 (.A(tie_lo_T8Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y35__R1_BUF_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R1_INV_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R2_INV_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y35__R2_INV_1 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y35__R3_BUF_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y36__R0_BUF_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R0_INV_0 (.A(tie_lo_T8Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y36__R1_BUF_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R1_INV_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R2_INV_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y36__R2_INV_1 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y36__R3_BUF_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y37__R0_BUF_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R0_INV_0 (.A(tie_lo_T8Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y37__R1_BUF_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R1_INV_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R2_INV_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y37__R2_INV_1 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y37__R3_BUF_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y38__R0_BUF_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R0_INV_0 (.A(tie_lo_T8Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y38__R1_BUF_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R1_INV_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R2_INV_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y38__R2_INV_1 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y38__R3_BUF_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y39__R0_BUF_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R0_INV_0 (.A(tie_lo_T8Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y39__R1_BUF_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R1_INV_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R2_INV_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y39__R2_INV_1 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y39__R3_BUF_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y3__R0_BUF_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R0_INV_0 (.A(tie_lo_T8Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y3__R1_BUF_0 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R1_INV_0 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R2_INV_0 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y3__R2_INV_1 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y3__R3_BUF_0 (.A(tie_lo_T8Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y40__R0_BUF_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R0_INV_0 (.A(tie_lo_T8Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y40__R1_BUF_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R1_INV_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R2_INV_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y40__R2_INV_1 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y40__R3_BUF_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y41__R0_BUF_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R0_INV_0 (.A(tie_lo_T8Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y41__R1_BUF_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R1_INV_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R2_INV_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y41__R2_INV_1 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y41__R3_BUF_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y42__R0_BUF_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R0_INV_0 (.A(tie_lo_T8Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y42__R1_BUF_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R1_INV_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R2_INV_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y42__R2_INV_1 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y42__R3_BUF_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y43__R0_BUF_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R0_INV_0 (.A(tie_lo_T8Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y43__R1_BUF_0 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R1_INV_0 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R2_INV_0 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y43__R2_INV_1 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y43__R3_BUF_0 (.A(tie_lo_T8Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y44__R0_BUF_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R0_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y44__R1_BUF_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R1_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R2_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y44__R2_INV_1 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y44__R3_BUF_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y45__R0_BUF_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R0_INV_0 (.A(tie_lo_T8Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y45__R1_BUF_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R1_INV_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R2_INV_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y45__R2_INV_1 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y45__R3_BUF_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y46__R0_BUF_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R0_INV_0 (.A(tie_lo_T8Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y46__R1_BUF_0 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R1_INV_0 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R2_INV_0 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y46__R2_INV_1 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y46__R3_BUF_0 (.A(tie_lo_T8Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y47__R0_BUF_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R0_INV_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y47__R1_BUF_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R1_INV_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R2_INV_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y47__R2_INV_1 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y47__R3_BUF_0 (.A(tie_lo_T8Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y48__R0_BUF_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R0_INV_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y48__R1_BUF_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R1_INV_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R2_INV_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y48__R2_INV_1 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y48__R3_BUF_0 (.A(tie_lo_T8Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y49__R0_BUF_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R0_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y49__R1_BUF_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R1_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R2_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y49__R2_INV_1 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y49__R3_BUF_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y4__R0_BUF_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R0_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y4__R1_BUF_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R1_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R2_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y4__R2_INV_1 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y4__R3_BUF_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y50__R0_BUF_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R0_INV_0 (.A(tie_lo_T8Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y50__R1_BUF_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R1_INV_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R2_INV_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y50__R2_INV_1 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y50__R3_BUF_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y51__R0_BUF_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R0_INV_0 (.A(tie_lo_T8Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y51__R1_BUF_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R1_INV_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R2_INV_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y51__R2_INV_1 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y51__R3_BUF_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y52__R0_BUF_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R0_INV_0 (.A(tie_lo_T8Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y52__R1_BUF_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R1_INV_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R2_INV_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y52__R2_INV_1 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y52__R3_BUF_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y53__R0_BUF_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R0_INV_0 (.A(tie_lo_T8Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y53__R1_BUF_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R1_INV_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R2_INV_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y53__R2_INV_1 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y53__R3_BUF_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y54__R0_BUF_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R0_INV_0 (.A(tie_lo_T8Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y54__R1_BUF_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R1_INV_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R2_INV_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y54__R2_INV_1 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y54__R3_BUF_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y55__R0_BUF_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R0_INV_0 (.A(tie_lo_T8Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y55__R1_BUF_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R1_INV_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R2_INV_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y55__R2_INV_1 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y55__R3_BUF_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y56__R0_BUF_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R0_INV_0 (.A(tie_lo_T8Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y56__R1_BUF_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R1_INV_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R2_INV_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y56__R2_INV_1 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y56__R3_BUF_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y57__R0_BUF_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R0_INV_0 (.A(tie_lo_T8Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y57__R1_BUF_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R1_INV_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R2_INV_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y57__R2_INV_1 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y57__R3_BUF_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y58__R0_BUF_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R0_INV_0 (.A(tie_lo_T8Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y58__R1_BUF_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R1_INV_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R2_INV_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y58__R2_INV_1 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y58__R3_BUF_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y59__R0_BUF_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R0_INV_0 (.A(tie_lo_T8Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y59__R1_BUF_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R1_INV_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R2_INV_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y59__R2_INV_1 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y59__R3_BUF_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y5__R0_BUF_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R0_INV_0 (.A(tie_lo_T8Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y5__R1_BUF_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R1_INV_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R2_INV_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y5__R2_INV_1 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y5__R3_BUF_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y60__R0_BUF_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R0_INV_0 (.A(tie_lo_T8Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y60__R1_BUF_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R1_INV_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R2_INV_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y60__R2_INV_1 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y60__R3_BUF_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y61__R0_BUF_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R0_INV_0 (.A(tie_lo_T8Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y61__R1_BUF_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R1_INV_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R2_INV_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y61__R2_INV_1 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y61__R3_BUF_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y62__R0_BUF_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R0_INV_0 (.A(tie_lo_T8Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y62__R1_BUF_0 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R1_INV_0 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R2_INV_0 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y62__R2_INV_1 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y62__R3_BUF_0 (.A(tie_lo_T8Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y63__R0_BUF_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R0_INV_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y63__R1_BUF_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R1_INV_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R2_INV_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y63__R2_INV_1 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y63__R3_BUF_0 (.A(tie_lo_T8Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y64__R0_BUF_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R0_INV_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y64__R1_BUF_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R1_INV_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R2_INV_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y64__R2_INV_1 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y64__R3_BUF_0 (.A(tie_lo_T8Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y65__R0_BUF_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R0_INV_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y65__R1_BUF_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R1_INV_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R2_INV_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y65__R2_INV_1 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y65__R3_BUF_0 (.A(tie_lo_T8Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y66__R0_BUF_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R0_INV_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y66__R1_BUF_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R1_INV_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R2_INV_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y66__R2_INV_1 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y66__R3_BUF_0 (.A(tie_lo_T8Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y67__R0_BUF_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R0_INV_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y67__R1_BUF_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R1_INV_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R2_INV_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y67__R2_INV_1 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y67__R3_BUF_0 (.A(tie_lo_T8Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y68__R0_BUF_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R0_INV_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y68__R1_BUF_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R1_INV_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R2_INV_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y68__R2_INV_1 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y68__R3_BUF_0 (.A(tie_lo_T8Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y69__R0_BUF_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R0_INV_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y69__R1_BUF_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R1_INV_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R2_INV_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y69__R2_INV_1 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y69__R3_BUF_0 (.A(tie_lo_T8Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y6__R0_BUF_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R0_INV_0 (.A(tie_lo_T8Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y6__R1_BUF_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R1_INV_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R2_INV_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y6__R2_INV_1 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y6__R3_BUF_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y70__R0_BUF_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R0_INV_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y70__R1_BUF_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R1_INV_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R2_INV_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y70__R2_INV_1 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y70__R3_BUF_0 (.A(tie_lo_T8Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y71__R0_BUF_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R0_INV_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y71__R1_BUF_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R1_INV_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R2_INV_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y71__R2_INV_1 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y71__R3_BUF_0 (.A(tie_lo_T8Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y72__R0_BUF_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R0_INV_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y72__R1_BUF_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R1_INV_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R2_INV_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y72__R2_INV_1 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y72__R3_BUF_0 (.A(tie_lo_T8Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y73__R0_BUF_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R0_INV_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y73__R1_BUF_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R1_INV_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R2_INV_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y73__R2_INV_1 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y73__R3_BUF_0 (.A(tie_lo_T8Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y74__R0_BUF_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R0_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y74__R1_BUF_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R1_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R2_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y74__R2_INV_1 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y74__R3_BUF_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y75__R0_BUF_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R0_INV_0 (.A(tie_lo_T8Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y75__R1_BUF_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R1_INV_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R2_INV_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y75__R2_INV_1 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y75__R3_BUF_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y76__R0_BUF_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R0_INV_0 (.A(tie_lo_T8Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y76__R1_BUF_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R1_INV_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R2_INV_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y76__R2_INV_1 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y76__R3_BUF_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y77__R0_BUF_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R0_INV_0 (.A(tie_lo_T8Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y77__R1_BUF_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R1_INV_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R2_INV_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y77__R2_INV_1 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y77__R3_BUF_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y78__R0_BUF_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R0_INV_0 (.A(tie_lo_T8Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y78__R1_BUF_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R1_INV_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R2_INV_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y78__R2_INV_1 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y78__R3_BUF_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y79__R0_BUF_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R0_INV_0 (.A(tie_lo_T8Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y79__R1_BUF_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R1_INV_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R2_INV_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y79__R2_INV_1 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y79__R3_BUF_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y7__R0_BUF_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R0_INV_0 (.A(tie_lo_T8Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y7__R1_BUF_0 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R1_INV_0 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R2_INV_0 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y7__R2_INV_1 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y7__R3_BUF_0 (.A(tie_lo_T8Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y80__R0_BUF_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R0_INV_0 (.A(tie_lo_T8Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y80__R1_BUF_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R1_INV_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R2_INV_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y80__R2_INV_1 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y80__R3_BUF_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y81__R0_BUF_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R0_INV_0 (.A(tie_lo_T8Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y81__R1_BUF_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R1_INV_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R2_INV_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y81__R2_INV_1 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y81__R3_BUF_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y82__R0_BUF_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R0_INV_0 (.A(tie_lo_T8Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y82__R1_BUF_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R1_INV_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R2_INV_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y82__R2_INV_1 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y82__R3_BUF_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y83__R0_BUF_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R0_INV_0 (.A(tie_lo_T8Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y83__R1_BUF_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R1_INV_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R2_INV_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y83__R2_INV_1 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y83__R3_BUF_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y84__R0_BUF_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R0_INV_0 (.A(tie_lo_T8Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y84__R1_BUF_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R1_INV_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R2_INV_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y84__R2_INV_1 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y84__R3_BUF_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y85__R0_BUF_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R0_INV_0 (.A(tie_lo_T8Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y85__R1_BUF_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R1_INV_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R2_INV_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y85__R2_INV_1 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y85__R3_BUF_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y86__R0_BUF_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R0_INV_0 (.A(tie_lo_T8Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y86__R1_BUF_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R1_INV_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R2_INV_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y86__R2_INV_1 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y86__R3_BUF_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y87__R0_BUF_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R0_INV_0 (.A(tie_lo_T8Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y87__R1_BUF_0 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R1_INV_0 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R2_INV_0 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y87__R2_INV_1 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y87__R3_BUF_0 (.A(tie_lo_T8Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y88__R0_BUF_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R0_INV_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y88__R1_BUF_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R1_INV_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R2_INV_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y88__R2_INV_1 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y88__R3_BUF_0 (.A(tie_lo_T8Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y89__R0_BUF_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R0_INV_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y89__R1_BUF_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R1_INV_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R2_INV_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y89__R2_INV_1 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y89__R3_BUF_0 (.A(tie_lo_T8Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y8__R0_BUF_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R0_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y8__R1_BUF_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R1_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R2_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y8__R2_INV_1 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y8__R3_BUF_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y9__R0_BUF_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R0_INV_0 (.A(tie_lo_T8Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y9__R1_BUF_0 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R1_INV_0 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T8Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R2_INV_0 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T8Y9__R2_INV_1 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T8Y9__R3_BUF_0 (.A(tie_lo_T8Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y0__R0_BUF_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R0_INV_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y0__R1_BUF_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R1_INV_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y0__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R2_INV_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y0__R2_INV_1 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y0__R3_BUF_0 (.A(tie_lo_T9Y0__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y10__R0_BUF_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R0_INV_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y10__R1_BUF_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R1_INV_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y10__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R2_INV_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y10__R2_INV_1 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y10__R3_BUF_0 (.A(tie_lo_T9Y10__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y11__R0_BUF_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R0_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y11__R1_BUF_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R1_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y11__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R2_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y11__R2_INV_1 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y11__R3_BUF_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y12__R0_BUF_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R0_INV_0 (.A(tie_lo_T9Y11__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y12__R1_BUF_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R1_INV_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y12__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R2_INV_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y12__R2_INV_1 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y12__R3_BUF_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y13__R0_BUF_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R0_INV_0 (.A(tie_lo_T9Y12__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y13__R1_BUF_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R1_INV_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y13__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R2_INV_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y13__R2_INV_1 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y13__R3_BUF_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y14__R0_BUF_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R0_INV_0 (.A(tie_lo_T9Y13__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y14__R1_BUF_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R1_INV_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y14__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R2_INV_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y14__R2_INV_1 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y14__R3_BUF_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y15__R0_BUF_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R0_INV_0 (.A(tie_lo_T9Y14__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y15__R1_BUF_0 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R1_INV_0 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y15__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R2_INV_0 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y15__R2_INV_1 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y15__R3_BUF_0 (.A(tie_lo_T9Y15__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y16__R0_BUF_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R0_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y16__R1_BUF_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R1_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y16__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R2_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y16__R2_INV_1 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y16__R3_BUF_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y17__R0_BUF_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R0_INV_0 (.A(tie_lo_T9Y16__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y17__R1_BUF_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R1_INV_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y17__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R2_INV_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y17__R2_INV_1 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y17__R3_BUF_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y18__R0_BUF_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R0_INV_0 (.A(tie_lo_T9Y17__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y18__R1_BUF_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R1_INV_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y18__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R2_INV_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y18__R2_INV_1 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y18__R3_BUF_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y19__R0_BUF_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R0_INV_0 (.A(tie_lo_T9Y18__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y19__R1_BUF_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R1_INV_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y19__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R2_INV_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y19__R2_INV_1 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y19__R3_BUF_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y1__R0_BUF_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R0_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y1__R1_BUF_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R1_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y1__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R2_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y1__R2_INV_1 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y1__R3_BUF_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y20__R0_BUF_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R0_INV_0 (.A(tie_lo_T9Y19__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y20__R1_BUF_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R1_INV_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y20__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R2_INV_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y20__R2_INV_1 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y20__R3_BUF_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y21__R0_BUF_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R0_INV_0 (.A(tie_lo_T9Y20__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y21__R1_BUF_0 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R1_INV_0 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y21__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R2_INV_0 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y21__R2_INV_1 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y21__R3_BUF_0 (.A(tie_lo_T9Y21__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y22__R0_BUF_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R0_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y22__R1_BUF_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R1_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y22__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R2_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y22__R2_INV_1 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y22__R3_BUF_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y23__R0_BUF_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R0_INV_0 (.A(tie_lo_T9Y22__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y23__R1_BUF_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R1_INV_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y23__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R2_INV_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y23__R2_INV_1 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y23__R3_BUF_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y24__R0_BUF_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R0_INV_0 (.A(tie_lo_T9Y23__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y24__R1_BUF_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R1_INV_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y24__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R2_INV_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y24__R2_INV_1 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y24__R3_BUF_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y25__R0_BUF_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R0_INV_0 (.A(tie_lo_T9Y24__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y25__R1_BUF_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R1_INV_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y25__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R2_INV_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y25__R2_INV_1 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y25__R3_BUF_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y26__R0_BUF_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R0_INV_0 (.A(tie_lo_T9Y25__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y26__R1_BUF_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R1_INV_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y26__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R2_INV_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y26__R2_INV_1 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y26__R3_BUF_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y27__R0_BUF_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R0_INV_0 (.A(tie_lo_T9Y26__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y27__R1_BUF_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R1_INV_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y27__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R2_INV_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y27__R2_INV_1 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y27__R3_BUF_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y28__R0_BUF_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R0_INV_0 (.A(tie_lo_T9Y27__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y28__R1_BUF_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R1_INV_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y28__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R2_INV_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y28__R2_INV_1 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y28__R3_BUF_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y29__R0_BUF_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R0_INV_0 (.A(tie_lo_T9Y28__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y29__R1_BUF_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R1_INV_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y29__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R2_INV_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y29__R2_INV_1 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y29__R3_BUF_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y2__R0_BUF_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R0_INV_0 (.A(tie_lo_T9Y1__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y2__R1_BUF_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R1_INV_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y2__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R2_INV_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y2__R2_INV_1 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y2__R3_BUF_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y30__R0_BUF_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R0_INV_0 (.A(tie_lo_T9Y29__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y30__R1_BUF_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R1_INV_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y30__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R2_INV_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y30__R2_INV_1 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y30__R3_BUF_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y31__R0_BUF_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R0_INV_0 (.A(tie_lo_T9Y30__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y31__R1_BUF_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R1_INV_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y31__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R2_INV_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y31__R2_INV_1 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y31__R3_BUF_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y32__R0_BUF_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R0_INV_0 (.A(tie_lo_T9Y31__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y32__R1_BUF_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R1_INV_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y32__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R2_INV_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y32__R2_INV_1 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y32__R3_BUF_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y33__R0_BUF_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R0_INV_0 (.A(tie_lo_T9Y32__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y33__R1_BUF_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R1_INV_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y33__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R2_INV_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y33__R2_INV_1 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y33__R3_BUF_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y34__R0_BUF_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R0_INV_0 (.A(tie_lo_T9Y33__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y34__R1_BUF_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R1_INV_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y34__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R2_INV_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y34__R2_INV_1 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y34__R3_BUF_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y35__R0_BUF_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R0_INV_0 (.A(tie_lo_T9Y34__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y35__R1_BUF_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R1_INV_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y35__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R2_INV_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y35__R2_INV_1 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y35__R3_BUF_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y36__R0_BUF_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R0_INV_0 (.A(tie_lo_T9Y35__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y36__R1_BUF_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R1_INV_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y36__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R2_INV_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y36__R2_INV_1 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y36__R3_BUF_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y37__R0_BUF_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R0_INV_0 (.A(tie_lo_T9Y36__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y37__R1_BUF_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R1_INV_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y37__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R2_INV_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y37__R2_INV_1 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y37__R3_BUF_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y38__R0_BUF_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R0_INV_0 (.A(tie_lo_T9Y37__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y38__R1_BUF_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R1_INV_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y38__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R2_INV_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y38__R2_INV_1 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y38__R3_BUF_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y39__R0_BUF_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R0_INV_0 (.A(tie_lo_T9Y38__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y39__R1_BUF_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R1_INV_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y39__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R2_INV_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y39__R2_INV_1 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y39__R3_BUF_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y3__R0_BUF_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R0_INV_0 (.A(tie_lo_T9Y2__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y3__R1_BUF_0 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R1_INV_0 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y3__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R2_INV_0 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y3__R2_INV_1 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y3__R3_BUF_0 (.A(tie_lo_T9Y3__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y40__R0_BUF_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R0_INV_0 (.A(tie_lo_T9Y39__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y40__R1_BUF_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R1_INV_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y40__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R2_INV_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y40__R2_INV_1 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y40__R3_BUF_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y41__R0_BUF_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R0_INV_0 (.A(tie_lo_T9Y40__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y41__R1_BUF_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R1_INV_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y41__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R2_INV_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y41__R2_INV_1 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y41__R3_BUF_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y42__R0_BUF_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R0_INV_0 (.A(tie_lo_T9Y41__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y42__R1_BUF_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R1_INV_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y42__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R2_INV_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y42__R2_INV_1 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y42__R3_BUF_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y43__R0_BUF_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R0_INV_0 (.A(tie_lo_T9Y42__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y43__R1_BUF_0 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R1_INV_0 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y43__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R2_INV_0 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y43__R2_INV_1 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y43__R3_BUF_0 (.A(tie_lo_T9Y43__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y44__R0_BUF_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R0_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y44__R1_BUF_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R1_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y44__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R2_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y44__R2_INV_1 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y44__R3_BUF_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y45__R0_BUF_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R0_INV_0 (.A(tie_lo_T9Y44__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y45__R1_BUF_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R1_INV_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y45__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R2_INV_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y45__R2_INV_1 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y45__R3_BUF_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y46__R0_BUF_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R0_INV_0 (.A(tie_lo_T9Y45__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y46__R1_BUF_0 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R1_INV_0 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y46__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R2_INV_0 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y46__R2_INV_1 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y46__R3_BUF_0 (.A(tie_lo_T9Y46__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y47__R0_BUF_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R0_INV_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y47__R1_BUF_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R1_INV_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y47__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R2_INV_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y47__R2_INV_1 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y47__R3_BUF_0 (.A(tie_lo_T9Y47__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y48__R0_BUF_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R0_INV_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y48__R1_BUF_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R1_INV_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y48__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R2_INV_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y48__R2_INV_1 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y48__R3_BUF_0 (.A(tie_lo_T9Y48__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y49__R0_BUF_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R0_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y49__R1_BUF_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R1_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y49__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R2_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y49__R2_INV_1 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y49__R3_BUF_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y4__R0_BUF_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R0_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y4__R1_BUF_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R1_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y4__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R2_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y4__R2_INV_1 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y4__R3_BUF_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y50__R0_BUF_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R0_INV_0 (.A(tie_lo_T9Y49__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y50__R1_BUF_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R1_INV_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y50__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R2_INV_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y50__R2_INV_1 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y50__R3_BUF_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y51__R0_BUF_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R0_INV_0 (.A(tie_lo_T9Y50__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y51__R1_BUF_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R1_INV_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y51__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R2_INV_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y51__R2_INV_1 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y51__R3_BUF_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y52__R0_BUF_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R0_INV_0 (.A(tie_lo_T9Y51__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y52__R1_BUF_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R1_INV_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y52__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R2_INV_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y52__R2_INV_1 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y52__R3_BUF_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y53__R0_BUF_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R0_INV_0 (.A(tie_lo_T9Y52__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y53__R1_BUF_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R1_INV_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y53__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R2_INV_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y53__R2_INV_1 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y53__R3_BUF_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y54__R0_BUF_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R0_INV_0 (.A(tie_lo_T9Y53__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y54__R1_BUF_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R1_INV_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y54__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R2_INV_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y54__R2_INV_1 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y54__R3_BUF_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y55__R0_BUF_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R0_INV_0 (.A(tie_lo_T9Y54__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y55__R1_BUF_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R1_INV_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y55__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R2_INV_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y55__R2_INV_1 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y55__R3_BUF_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y56__R0_BUF_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R0_INV_0 (.A(tie_lo_T9Y55__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y56__R1_BUF_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R1_INV_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y56__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R2_INV_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y56__R2_INV_1 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y56__R3_BUF_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y57__R0_BUF_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R0_INV_0 (.A(tie_lo_T9Y56__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y57__R1_BUF_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R1_INV_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y57__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R2_INV_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y57__R2_INV_1 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y57__R3_BUF_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y58__R0_BUF_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R0_INV_0 (.A(tie_lo_T9Y57__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y58__R1_BUF_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R1_INV_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y58__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R2_INV_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y58__R2_INV_1 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y58__R3_BUF_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y59__R0_BUF_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R0_INV_0 (.A(tie_lo_T9Y58__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y59__R1_BUF_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R1_INV_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y59__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R2_INV_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y59__R2_INV_1 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y59__R3_BUF_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y5__R0_BUF_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R0_INV_0 (.A(tie_lo_T9Y4__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y5__R1_BUF_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R1_INV_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y5__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R2_INV_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y5__R2_INV_1 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y5__R3_BUF_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y60__R0_BUF_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R0_INV_0 (.A(tie_lo_T9Y59__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y60__R1_BUF_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R1_INV_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y60__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R2_INV_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y60__R2_INV_1 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y60__R3_BUF_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y61__R0_BUF_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R0_INV_0 (.A(tie_lo_T9Y60__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y61__R1_BUF_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R1_INV_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y61__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R2_INV_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y61__R2_INV_1 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y61__R3_BUF_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y62__R0_BUF_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R0_INV_0 (.A(tie_lo_T9Y61__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y62__R1_BUF_0 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R1_INV_0 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y62__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R2_INV_0 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y62__R2_INV_1 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y62__R3_BUF_0 (.A(tie_lo_T9Y62__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y63__R0_BUF_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R0_INV_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y63__R1_BUF_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R1_INV_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y63__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R2_INV_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y63__R2_INV_1 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y63__R3_BUF_0 (.A(tie_lo_T9Y63__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y64__R0_BUF_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R0_INV_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y64__R1_BUF_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R1_INV_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y64__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R2_INV_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y64__R2_INV_1 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y64__R3_BUF_0 (.A(tie_lo_T9Y64__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y65__R0_BUF_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R0_INV_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y65__R1_BUF_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R1_INV_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y65__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R2_INV_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y65__R2_INV_1 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y65__R3_BUF_0 (.A(tie_lo_T9Y65__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y66__R0_BUF_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R0_INV_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y66__R1_BUF_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R1_INV_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y66__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R2_INV_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y66__R2_INV_1 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y66__R3_BUF_0 (.A(tie_lo_T9Y66__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y67__R0_BUF_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R0_INV_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y67__R1_BUF_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R1_INV_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y67__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R2_INV_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y67__R2_INV_1 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y67__R3_BUF_0 (.A(tie_lo_T9Y67__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y68__R0_BUF_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R0_INV_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y68__R1_BUF_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R1_INV_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y68__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R2_INV_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y68__R2_INV_1 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y68__R3_BUF_0 (.A(tie_lo_T9Y68__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y69__R0_BUF_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R0_INV_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y69__R1_BUF_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R1_INV_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y69__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R2_INV_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y69__R2_INV_1 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y69__R3_BUF_0 (.A(tie_lo_T9Y69__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y6__R0_BUF_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R0_INV_0 (.A(tie_lo_T9Y5__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y6__R1_BUF_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R1_INV_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y6__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R2_INV_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y6__R2_INV_1 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y6__R3_BUF_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y70__R0_BUF_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R0_INV_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y70__R1_BUF_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R1_INV_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y70__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R2_INV_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y70__R2_INV_1 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y70__R3_BUF_0 (.A(tie_lo_T9Y70__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y71__R0_BUF_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R0_INV_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y71__R1_BUF_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R1_INV_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y71__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R2_INV_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y71__R2_INV_1 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y71__R3_BUF_0 (.A(tie_lo_T9Y71__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y72__R0_BUF_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R0_INV_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y72__R1_BUF_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R1_INV_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y72__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R2_INV_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y72__R2_INV_1 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y72__R3_BUF_0 (.A(tie_lo_T9Y72__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y73__R0_BUF_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R0_INV_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y73__R1_BUF_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R1_INV_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y73__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R2_INV_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y73__R2_INV_1 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y73__R3_BUF_0 (.A(tie_lo_T9Y73__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y74__R0_BUF_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R0_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y74__R1_BUF_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R1_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y74__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R2_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y74__R2_INV_1 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y74__R3_BUF_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y75__R0_BUF_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R0_INV_0 (.A(tie_lo_T9Y74__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y75__R1_BUF_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R1_INV_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y75__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R2_INV_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y75__R2_INV_1 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y75__R3_BUF_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y76__R0_BUF_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R0_INV_0 (.A(tie_lo_T9Y75__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y76__R1_BUF_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R1_INV_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y76__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R2_INV_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y76__R2_INV_1 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y76__R3_BUF_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y77__R0_BUF_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R0_INV_0 (.A(tie_lo_T9Y76__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y77__R1_BUF_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R1_INV_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y77__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R2_INV_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y77__R2_INV_1 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y77__R3_BUF_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y78__R0_BUF_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R0_INV_0 (.A(tie_lo_T9Y77__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y78__R1_BUF_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R1_INV_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y78__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R2_INV_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y78__R2_INV_1 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y78__R3_BUF_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y79__R0_BUF_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R0_INV_0 (.A(tie_lo_T9Y78__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y79__R1_BUF_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R1_INV_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y79__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R2_INV_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y79__R2_INV_1 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y79__R3_BUF_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y7__R0_BUF_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R0_INV_0 (.A(tie_lo_T9Y6__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y7__R1_BUF_0 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R1_INV_0 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y7__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R2_INV_0 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y7__R2_INV_1 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y7__R3_BUF_0 (.A(tie_lo_T9Y7__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y80__R0_BUF_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R0_INV_0 (.A(tie_lo_T9Y79__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y80__R1_BUF_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R1_INV_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y80__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R2_INV_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y80__R2_INV_1 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y80__R3_BUF_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y81__R0_BUF_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R0_INV_0 (.A(tie_lo_T9Y80__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y81__R1_BUF_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R1_INV_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y81__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R2_INV_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y81__R2_INV_1 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y81__R3_BUF_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y82__R0_BUF_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R0_INV_0 (.A(tie_lo_T9Y81__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y82__R1_BUF_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R1_INV_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y82__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R2_INV_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y82__R2_INV_1 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y82__R3_BUF_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y83__R0_BUF_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R0_INV_0 (.A(tie_lo_T9Y82__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y83__R1_BUF_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R1_INV_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y83__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R2_INV_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y83__R2_INV_1 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y83__R3_BUF_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y84__R0_BUF_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R0_INV_0 (.A(tie_lo_T9Y83__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y84__R1_BUF_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R1_INV_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y84__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R2_INV_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y84__R2_INV_1 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y84__R3_BUF_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y85__R0_BUF_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R0_INV_0 (.A(tie_lo_T9Y84__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y85__R1_BUF_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R1_INV_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y85__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R2_INV_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y85__R2_INV_1 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y85__R3_BUF_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y86__R0_BUF_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R0_INV_0 (.A(tie_lo_T9Y85__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y86__R1_BUF_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R1_INV_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y86__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R2_INV_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y86__R2_INV_1 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y86__R3_BUF_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y87__R0_BUF_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R0_INV_0 (.A(tie_lo_T9Y86__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y87__R1_BUF_0 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R1_INV_0 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y87__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R2_INV_0 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y87__R2_INV_1 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y87__R3_BUF_0 (.A(tie_lo_T9Y87__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y88__R0_BUF_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R0_INV_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y88__R1_BUF_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R1_INV_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y88__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R2_INV_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y88__R2_INV_1 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y88__R3_BUF_0 (.A(tie_lo_T9Y88__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y89__R0_BUF_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R0_INV_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y89__R1_BUF_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R1_INV_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y89__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R2_INV_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y89__R2_INV_1 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y89__R3_BUF_0 (.A(tie_lo_T9Y89__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y8__R0_BUF_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R0_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y8__R1_BUF_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R1_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y8__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R2_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y8__R2_INV_1 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y8__R3_BUF_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y9__R0_BUF_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R0_INV_0 (.A(tie_lo_T9Y8__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y9__R1_BUF_0 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R1_INV_0 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__conb_1 T9Y9__R2_CONB_0 (.HI(vdd_unused), .LO(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R2_INV_0 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkinv_2 T9Y9__R2_INV_1 (.A(tie_lo_T9Y9__R2_CONB_0));
  sky130_fd_sc_hd__clkbuf_4 T9Y9__R3_BUF_0 (.A(tie_lo_T9Y9__R2_CONB_0));

endmodule
