module sasic_top (
  clk,
  rst_n,
  in_0,
  in_1,
  in_2,
  in_3,
  in_4,
  in_5,
  in_6,
  in_7,
  in_8,
  in_9,
  in_10,
  in_11,
  in_12,
  in_13,
  in_14,
  in_15,
  in_16,
  in_17,
  in_18,
  in_19,
  in_20,
  in_21,
  in_22,
  in_23,
  in_24,
  in_25,
  in_26,
  in_27,
  in_28,
  in_29,
  in_30,
  in_31,
  in_32,
  in_33,
  in_34,
  in_35,
  in_36,
  in_37,
  in_38,
  in_39,
  oeb_0,
  oeb_1,
  oeb_2,
  oeb_3,
  oeb_4,
  oeb_5,
  oeb_6,
  oeb_7,
  oeb_8,
  oeb_9,
  oeb_10,
  oeb_11,
  oeb_12,
  oeb_13,
  oeb_14,
  oeb_15,
  oeb_16,
  oeb_17,
  oeb_18,
  oeb_19,
  oeb_20,
  oeb_21,
  oeb_22,
  oeb_23,
  oeb_24,
  oeb_25,
  oeb_26,
  oeb_27,
  oeb_28,
  oeb_29,
  oeb_30,
  oeb_31,
  oeb_32,
  oeb_33,
  oeb_34,
  oeb_35,
  oeb_36,
  oeb_37,
  oeb_38,
  oeb_39,
  out_0,
  out_1,
  out_2,
  out_3,
  out_4,
  out_5,
  out_6,
  out_7,
  out_8,
  out_9,
  out_10,
  out_11,
  out_12,
  out_13,
  out_14,
  out_15,
  out_16,
  out_17,
  out_18,
  out_19,
  out_20,
  out_21,
  out_22,
  out_23,
  out_24,
  out_25,
  out_26,
  out_27,
  out_28,
  out_29,
  out_30,
  out_31,
  out_32,
  out_33,
  out_34,
  out_35,
  out_36,
  out_37,
  out_38,
  out_39
);

  input clk;
  input rst_n;
  input in_0;
  input in_1;
  input in_2;
  input in_3;
  input in_4;
  input in_5;
  input in_6;
  input in_7;
  input in_8;
  input in_9;
  input in_10;
  input in_11;
  input in_12;
  input in_13;
  input in_14;
  input in_15;
  input in_16;
  input in_17;
  input in_18;
  input in_19;
  input in_20;
  input in_21;
  input in_22;
  input in_23;
  input in_24;
  input in_25;
  input in_26;
  input in_27;
  input in_28;
  input in_29;
  input in_30;
  input in_31;
  input in_32;
  input in_33;
  input in_34;
  input in_35;
  input in_36;
  input in_37;
  input in_38;
  input in_39;
  output oeb_0;
  output oeb_1;
  output oeb_2;
  output oeb_3;
  output oeb_4;
  output oeb_5;
  output oeb_6;
  output oeb_7;
  output oeb_8;
  output oeb_9;
  output oeb_10;
  output oeb_11;
  output oeb_12;
  output oeb_13;
  output oeb_14;
  output oeb_15;
  output oeb_16;
  output oeb_17;
  output oeb_18;
  output oeb_19;
  output oeb_20;
  output oeb_21;
  output oeb_22;
  output oeb_23;
  output oeb_24;
  output oeb_25;
  output oeb_26;
  output oeb_27;
  output oeb_28;
  output oeb_29;
  output oeb_30;
  output oeb_31;
  output oeb_32;
  output oeb_33;
  output oeb_34;
  output oeb_35;
  output oeb_36;
  output oeb_37;
  output oeb_38;
  output oeb_39;
  output out_0;
  output out_1;
  output out_2;
  output out_3;
  output out_4;
  output out_5;
  output out_6;
  output out_7;
  output out_8;
  output out_9;
  output out_10;
  output out_11;
  output out_12;
  output out_13;
  output out_14;
  output out_15;
  output out_16;
  output out_17;
  output out_18;
  output out_19;
  output out_20;
  output out_21;
  output out_22;
  output out_23;
  output out_24;
  output out_25;
  output out_26;
  output out_27;
  output out_28;
  output out_29;
  output out_30;
  output out_31;
  output out_32;
  output out_33;
  output out_34;
  output out_35;
  output out_36;
  output out_37;
  output out_38;
  output out_39;

  // Internal nets
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9110 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9120 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9132 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9134 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9136 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9138 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9140 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9142 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9174 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9180 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9182 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9184 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9210 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9226 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9228 ;
  wire \$abc$9276$auto$dfflibmap.cc:532:dfflibmap$9264 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8819 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8821 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8823 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8825 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8827 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8829 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8831 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8833 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8835 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8837 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8839 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8841 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8843 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8845 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8847 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8849 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8851 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8853 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8855 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8857 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8859 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8861 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8863 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8865 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8867 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8869 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8871 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8873 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8875 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8877 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8879 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8881 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8883 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8887 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8889 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8891 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8893 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8895 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8897 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8899 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8901 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8903 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8905 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8907 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8909 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8911 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8913 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8915 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8917 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8921 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8923 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8925 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8927 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8929 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8931 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8933 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8935 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8937 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8939 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8941 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8943 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8945 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8947 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8949 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8951 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8953 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8955 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8957 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8959 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8961 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8963 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8965 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8969 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8971 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8973 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8975 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8979 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8981 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8983 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8987 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8989 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8991 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8993 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8995 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8997 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$8999 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9001 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9003 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9005 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9007 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9009 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9011 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9013 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9015 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9017 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9019 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9021 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9023 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9025 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9027 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9029 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9031 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9033 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9035 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9037 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9039 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9041 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9043 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9045 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9047 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9049 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9051 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9053 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9057 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9061 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9065 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9069 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9073 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9077 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9081 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9085 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9087 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9089 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9091 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9093 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9095 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9097 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9099 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9101 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9103 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9105 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9107 ;
  wire \$abc$9276$auto$rtlil.cc:3205:MuxGate$9109 ;
  wire \$abc$9276$flatten \CPU.\$0 \adj_bcd[0:0];
  wire \$abc$9276$new_n1000 ;
  wire \$abc$9276$new_n1001 ;
  wire \$abc$9276$new_n1002 ;
  wire \$abc$9276$new_n1003 ;
  wire \$abc$9276$new_n1004 ;
  wire \$abc$9276$new_n1005 ;
  wire \$abc$9276$new_n1006 ;
  wire \$abc$9276$new_n1007 ;
  wire \$abc$9276$new_n1008 ;
  wire \$abc$9276$new_n1009 ;
  wire \$abc$9276$new_n1010 ;
  wire \$abc$9276$new_n1011 ;
  wire \$abc$9276$new_n1012 ;
  wire \$abc$9276$new_n1013 ;
  wire \$abc$9276$new_n1014 ;
  wire \$abc$9276$new_n1015 ;
  wire \$abc$9276$new_n1016 ;
  wire \$abc$9276$new_n1017 ;
  wire \$abc$9276$new_n1018 ;
  wire \$abc$9276$new_n1019 ;
  wire \$abc$9276$new_n1020 ;
  wire \$abc$9276$new_n1021 ;
  wire \$abc$9276$new_n1022 ;
  wire \$abc$9276$new_n1023 ;
  wire \$abc$9276$new_n1024 ;
  wire \$abc$9276$new_n1025 ;
  wire \$abc$9276$new_n1026 ;
  wire \$abc$9276$new_n1027 ;
  wire \$abc$9276$new_n1028 ;
  wire \$abc$9276$new_n1029 ;
  wire \$abc$9276$new_n1030 ;
  wire \$abc$9276$new_n1031 ;
  wire \$abc$9276$new_n1032 ;
  wire \$abc$9276$new_n1033 ;
  wire \$abc$9276$new_n1034 ;
  wire \$abc$9276$new_n1035 ;
  wire \$abc$9276$new_n1036 ;
  wire \$abc$9276$new_n1037 ;
  wire \$abc$9276$new_n1039 ;
  wire \$abc$9276$new_n1040 ;
  wire \$abc$9276$new_n1041 ;
  wire \$abc$9276$new_n1042 ;
  wire \$abc$9276$new_n1043 ;
  wire \$abc$9276$new_n1044 ;
  wire \$abc$9276$new_n1045 ;
  wire \$abc$9276$new_n1046 ;
  wire \$abc$9276$new_n1047 ;
  wire \$abc$9276$new_n1048 ;
  wire \$abc$9276$new_n1049 ;
  wire \$abc$9276$new_n1050 ;
  wire \$abc$9276$new_n1051 ;
  wire \$abc$9276$new_n1052 ;
  wire \$abc$9276$new_n1053 ;
  wire \$abc$9276$new_n1054 ;
  wire \$abc$9276$new_n1055 ;
  wire \$abc$9276$new_n1056 ;
  wire \$abc$9276$new_n1058 ;
  wire \$abc$9276$new_n1059 ;
  wire \$abc$9276$new_n1060 ;
  wire \$abc$9276$new_n1061 ;
  wire \$abc$9276$new_n1062 ;
  wire \$abc$9276$new_n1063 ;
  wire \$abc$9276$new_n1064 ;
  wire \$abc$9276$new_n1065 ;
  wire \$abc$9276$new_n1066 ;
  wire \$abc$9276$new_n1067 ;
  wire \$abc$9276$new_n1068 ;
  wire \$abc$9276$new_n1069 ;
  wire \$abc$9276$new_n1070 ;
  wire \$abc$9276$new_n1071 ;
  wire \$abc$9276$new_n1072 ;
  wire \$abc$9276$new_n1073 ;
  wire \$abc$9276$new_n1074 ;
  wire \$abc$9276$new_n1075 ;
  wire \$abc$9276$new_n1076 ;
  wire \$abc$9276$new_n1077 ;
  wire \$abc$9276$new_n1078 ;
  wire \$abc$9276$new_n1079 ;
  wire \$abc$9276$new_n1081 ;
  wire \$abc$9276$new_n1082 ;
  wire \$abc$9276$new_n1083 ;
  wire \$abc$9276$new_n1084 ;
  wire \$abc$9276$new_n1085 ;
  wire \$abc$9276$new_n1086 ;
  wire \$abc$9276$new_n1087 ;
  wire \$abc$9276$new_n1088 ;
  wire \$abc$9276$new_n1089 ;
  wire \$abc$9276$new_n1090 ;
  wire \$abc$9276$new_n1091 ;
  wire \$abc$9276$new_n1092 ;
  wire \$abc$9276$new_n1093 ;
  wire \$abc$9276$new_n1094 ;
  wire \$abc$9276$new_n1095 ;
  wire \$abc$9276$new_n1096 ;
  wire \$abc$9276$new_n1098 ;
  wire \$abc$9276$new_n1099 ;
  wire \$abc$9276$new_n1100 ;
  wire \$abc$9276$new_n1101 ;
  wire \$abc$9276$new_n1102 ;
  wire \$abc$9276$new_n1103 ;
  wire \$abc$9276$new_n1104 ;
  wire \$abc$9276$new_n1105 ;
  wire \$abc$9276$new_n1106 ;
  wire \$abc$9276$new_n1107 ;
  wire \$abc$9276$new_n1108 ;
  wire \$abc$9276$new_n1109 ;
  wire \$abc$9276$new_n1110 ;
  wire \$abc$9276$new_n1111 ;
  wire \$abc$9276$new_n1112 ;
  wire \$abc$9276$new_n1113 ;
  wire \$abc$9276$new_n1115 ;
  wire \$abc$9276$new_n1116 ;
  wire \$abc$9276$new_n1117 ;
  wire \$abc$9276$new_n1118 ;
  wire \$abc$9276$new_n1119 ;
  wire \$abc$9276$new_n1120 ;
  wire \$abc$9276$new_n1121 ;
  wire \$abc$9276$new_n1122 ;
  wire \$abc$9276$new_n1123 ;
  wire \$abc$9276$new_n1124 ;
  wire \$abc$9276$new_n1125 ;
  wire \$abc$9276$new_n1126 ;
  wire \$abc$9276$new_n1127 ;
  wire \$abc$9276$new_n1128 ;
  wire \$abc$9276$new_n1129 ;
  wire \$abc$9276$new_n1130 ;
  wire \$abc$9276$new_n1131 ;
  wire \$abc$9276$new_n1133 ;
  wire \$abc$9276$new_n1134 ;
  wire \$abc$9276$new_n1135 ;
  wire \$abc$9276$new_n1136 ;
  wire \$abc$9276$new_n1137 ;
  wire \$abc$9276$new_n1138 ;
  wire \$abc$9276$new_n1139 ;
  wire \$abc$9276$new_n1140 ;
  wire \$abc$9276$new_n1141 ;
  wire \$abc$9276$new_n1142 ;
  wire \$abc$9276$new_n1143 ;
  wire \$abc$9276$new_n1144 ;
  wire \$abc$9276$new_n1145 ;
  wire \$abc$9276$new_n1146 ;
  wire \$abc$9276$new_n1147 ;
  wire \$abc$9276$new_n1148 ;
  wire \$abc$9276$new_n1150 ;
  wire \$abc$9276$new_n1151 ;
  wire \$abc$9276$new_n1152 ;
  wire \$abc$9276$new_n1153 ;
  wire \$abc$9276$new_n1154 ;
  wire \$abc$9276$new_n1155 ;
  wire \$abc$9276$new_n1156 ;
  wire \$abc$9276$new_n1157 ;
  wire \$abc$9276$new_n1158 ;
  wire \$abc$9276$new_n1159 ;
  wire \$abc$9276$new_n1160 ;
  wire \$abc$9276$new_n1161 ;
  wire \$abc$9276$new_n1162 ;
  wire \$abc$9276$new_n1163 ;
  wire \$abc$9276$new_n1164 ;
  wire \$abc$9276$new_n1165 ;
  wire \$abc$9276$new_n1167 ;
  wire \$abc$9276$new_n1168 ;
  wire \$abc$9276$new_n1169 ;
  wire \$abc$9276$new_n1170 ;
  wire \$abc$9276$new_n1171 ;
  wire \$abc$9276$new_n1172 ;
  wire \$abc$9276$new_n1173 ;
  wire \$abc$9276$new_n1174 ;
  wire \$abc$9276$new_n1175 ;
  wire \$abc$9276$new_n1176 ;
  wire \$abc$9276$new_n1177 ;
  wire \$abc$9276$new_n1178 ;
  wire \$abc$9276$new_n1179 ;
  wire \$abc$9276$new_n1180 ;
  wire \$abc$9276$new_n1181 ;
  wire \$abc$9276$new_n1182 ;
  wire \$abc$9276$new_n1183 ;
  wire \$abc$9276$new_n1184 ;
  wire \$abc$9276$new_n1185 ;
  wire \$abc$9276$new_n1187 ;
  wire \$abc$9276$new_n1188 ;
  wire \$abc$9276$new_n1189 ;
  wire \$abc$9276$new_n1190 ;
  wire \$abc$9276$new_n1191 ;
  wire \$abc$9276$new_n1192 ;
  wire \$abc$9276$new_n1193 ;
  wire \$abc$9276$new_n1194 ;
  wire \$abc$9276$new_n1195 ;
  wire \$abc$9276$new_n1196 ;
  wire \$abc$9276$new_n1197 ;
  wire \$abc$9276$new_n1198 ;
  wire \$abc$9276$new_n1199 ;
  wire \$abc$9276$new_n1200 ;
  wire \$abc$9276$new_n1201 ;
  wire \$abc$9276$new_n1202 ;
  wire \$abc$9276$new_n1203 ;
  wire \$abc$9276$new_n1204 ;
  wire \$abc$9276$new_n1206 ;
  wire \$abc$9276$new_n1207 ;
  wire \$abc$9276$new_n1208 ;
  wire \$abc$9276$new_n1209 ;
  wire \$abc$9276$new_n1210 ;
  wire \$abc$9276$new_n1211 ;
  wire \$abc$9276$new_n1212 ;
  wire \$abc$9276$new_n1213 ;
  wire \$abc$9276$new_n1214 ;
  wire \$abc$9276$new_n1215 ;
  wire \$abc$9276$new_n1216 ;
  wire \$abc$9276$new_n1217 ;
  wire \$abc$9276$new_n1218 ;
  wire \$abc$9276$new_n1219 ;
  wire \$abc$9276$new_n1220 ;
  wire \$abc$9276$new_n1221 ;
  wire \$abc$9276$new_n1222 ;
  wire \$abc$9276$new_n1223 ;
  wire \$abc$9276$new_n1224 ;
  wire \$abc$9276$new_n1226 ;
  wire \$abc$9276$new_n1227 ;
  wire \$abc$9276$new_n1228 ;
  wire \$abc$9276$new_n1229 ;
  wire \$abc$9276$new_n1230 ;
  wire \$abc$9276$new_n1231 ;
  wire \$abc$9276$new_n1232 ;
  wire \$abc$9276$new_n1233 ;
  wire \$abc$9276$new_n1234 ;
  wire \$abc$9276$new_n1235 ;
  wire \$abc$9276$new_n1236 ;
  wire \$abc$9276$new_n1237 ;
  wire \$abc$9276$new_n1238 ;
  wire \$abc$9276$new_n1239 ;
  wire \$abc$9276$new_n1240 ;
  wire \$abc$9276$new_n1241 ;
  wire \$abc$9276$new_n1242 ;
  wire \$abc$9276$new_n1243 ;
  wire \$abc$9276$new_n1245 ;
  wire \$abc$9276$new_n1246 ;
  wire \$abc$9276$new_n1247 ;
  wire \$abc$9276$new_n1248 ;
  wire \$abc$9276$new_n1249 ;
  wire \$abc$9276$new_n1250 ;
  wire \$abc$9276$new_n1251 ;
  wire \$abc$9276$new_n1252 ;
  wire \$abc$9276$new_n1253 ;
  wire \$abc$9276$new_n1254 ;
  wire \$abc$9276$new_n1255 ;
  wire \$abc$9276$new_n1256 ;
  wire \$abc$9276$new_n1257 ;
  wire \$abc$9276$new_n1258 ;
  wire \$abc$9276$new_n1259 ;
  wire \$abc$9276$new_n1260 ;
  wire \$abc$9276$new_n1261 ;
  wire \$abc$9276$new_n1262 ;
  wire \$abc$9276$new_n1263 ;
  wire \$abc$9276$new_n1264 ;
  wire \$abc$9276$new_n1266 ;
  wire \$abc$9276$new_n1267 ;
  wire \$abc$9276$new_n1268 ;
  wire \$abc$9276$new_n1269 ;
  wire \$abc$9276$new_n1270 ;
  wire \$abc$9276$new_n1271 ;
  wire \$abc$9276$new_n1272 ;
  wire \$abc$9276$new_n1273 ;
  wire \$abc$9276$new_n1274 ;
  wire \$abc$9276$new_n1275 ;
  wire \$abc$9276$new_n1276 ;
  wire \$abc$9276$new_n1277 ;
  wire \$abc$9276$new_n1278 ;
  wire \$abc$9276$new_n1279 ;
  wire \$abc$9276$new_n1280 ;
  wire \$abc$9276$new_n1281 ;
  wire \$abc$9276$new_n1282 ;
  wire \$abc$9276$new_n1283 ;
  wire \$abc$9276$new_n1284 ;
  wire \$abc$9276$new_n1286 ;
  wire \$abc$9276$new_n1287 ;
  wire \$abc$9276$new_n1288 ;
  wire \$abc$9276$new_n1289 ;
  wire \$abc$9276$new_n1290 ;
  wire \$abc$9276$new_n1291 ;
  wire \$abc$9276$new_n1292 ;
  wire \$abc$9276$new_n1293 ;
  wire \$abc$9276$new_n1294 ;
  wire \$abc$9276$new_n1295 ;
  wire \$abc$9276$new_n1296 ;
  wire \$abc$9276$new_n1297 ;
  wire \$abc$9276$new_n1298 ;
  wire \$abc$9276$new_n1299 ;
  wire \$abc$9276$new_n1300 ;
  wire \$abc$9276$new_n1301 ;
  wire \$abc$9276$new_n1302 ;
  wire \$abc$9276$new_n1304 ;
  wire \$abc$9276$new_n1305 ;
  wire \$abc$9276$new_n1306 ;
  wire \$abc$9276$new_n1307 ;
  wire \$abc$9276$new_n1308 ;
  wire \$abc$9276$new_n1309 ;
  wire \$abc$9276$new_n1310 ;
  wire \$abc$9276$new_n1311 ;
  wire \$abc$9276$new_n1312 ;
  wire \$abc$9276$new_n1313 ;
  wire \$abc$9276$new_n1314 ;
  wire \$abc$9276$new_n1315 ;
  wire \$abc$9276$new_n1316 ;
  wire \$abc$9276$new_n1317 ;
  wire \$abc$9276$new_n1318 ;
  wire \$abc$9276$new_n1319 ;
  wire \$abc$9276$new_n1321 ;
  wire \$abc$9276$new_n1322 ;
  wire \$abc$9276$new_n1324 ;
  wire \$abc$9276$new_n1325 ;
  wire \$abc$9276$new_n1327 ;
  wire \$abc$9276$new_n1328 ;
  wire \$abc$9276$new_n1330 ;
  wire \$abc$9276$new_n1331 ;
  wire \$abc$9276$new_n1332 ;
  wire \$abc$9276$new_n1333 ;
  wire \$abc$9276$new_n1334 ;
  wire \$abc$9276$new_n1335 ;
  wire \$abc$9276$new_n1336 ;
  wire \$abc$9276$new_n1337 ;
  wire \$abc$9276$new_n1338 ;
  wire \$abc$9276$new_n1339 ;
  wire \$abc$9276$new_n1340 ;
  wire \$abc$9276$new_n1341 ;
  wire \$abc$9276$new_n1342 ;
  wire \$abc$9276$new_n1343 ;
  wire \$abc$9276$new_n1344 ;
  wire \$abc$9276$new_n1345 ;
  wire \$abc$9276$new_n1347 ;
  wire \$abc$9276$new_n1348 ;
  wire \$abc$9276$new_n1349 ;
  wire \$abc$9276$new_n1350 ;
  wire \$abc$9276$new_n1351 ;
  wire \$abc$9276$new_n1352 ;
  wire \$abc$9276$new_n1353 ;
  wire \$abc$9276$new_n1354 ;
  wire \$abc$9276$new_n1355 ;
  wire \$abc$9276$new_n1356 ;
  wire \$abc$9276$new_n1357 ;
  wire \$abc$9276$new_n1358 ;
  wire \$abc$9276$new_n1359 ;
  wire \$abc$9276$new_n1360 ;
  wire \$abc$9276$new_n1361 ;
  wire \$abc$9276$new_n1362 ;
  wire \$abc$9276$new_n1363 ;
  wire \$abc$9276$new_n1364 ;
  wire \$abc$9276$new_n1366 ;
  wire \$abc$9276$new_n1367 ;
  wire \$abc$9276$new_n1368 ;
  wire \$abc$9276$new_n1369 ;
  wire \$abc$9276$new_n1370 ;
  wire \$abc$9276$new_n1371 ;
  wire \$abc$9276$new_n1372 ;
  wire \$abc$9276$new_n1373 ;
  wire \$abc$9276$new_n1374 ;
  wire \$abc$9276$new_n1375 ;
  wire \$abc$9276$new_n1376 ;
  wire \$abc$9276$new_n1377 ;
  wire \$abc$9276$new_n1378 ;
  wire \$abc$9276$new_n1379 ;
  wire \$abc$9276$new_n1380 ;
  wire \$abc$9276$new_n1381 ;
  wire \$abc$9276$new_n1382 ;
  wire \$abc$9276$new_n1383 ;
  wire \$abc$9276$new_n1384 ;
  wire \$abc$9276$new_n1385 ;
  wire \$abc$9276$new_n1386 ;
  wire \$abc$9276$new_n1387 ;
  wire \$abc$9276$new_n1388 ;
  wire \$abc$9276$new_n1389 ;
  wire \$abc$9276$new_n1390 ;
  wire \$abc$9276$new_n1392 ;
  wire \$abc$9276$new_n1393 ;
  wire \$abc$9276$new_n1394 ;
  wire \$abc$9276$new_n1395 ;
  wire \$abc$9276$new_n1396 ;
  wire \$abc$9276$new_n1397 ;
  wire \$abc$9276$new_n1398 ;
  wire \$abc$9276$new_n1399 ;
  wire \$abc$9276$new_n1400 ;
  wire \$abc$9276$new_n1401 ;
  wire \$abc$9276$new_n1402 ;
  wire \$abc$9276$new_n1403 ;
  wire \$abc$9276$new_n1404 ;
  wire \$abc$9276$new_n1405 ;
  wire \$abc$9276$new_n1406 ;
  wire \$abc$9276$new_n1407 ;
  wire \$abc$9276$new_n1408 ;
  wire \$abc$9276$new_n1409 ;
  wire \$abc$9276$new_n1410 ;
  wire \$abc$9276$new_n1411 ;
  wire \$abc$9276$new_n1412 ;
  wire \$abc$9276$new_n1413 ;
  wire \$abc$9276$new_n1414 ;
  wire \$abc$9276$new_n1415 ;
  wire \$abc$9276$new_n1416 ;
  wire \$abc$9276$new_n1417 ;
  wire \$abc$9276$new_n1418 ;
  wire \$abc$9276$new_n1419 ;
  wire \$abc$9276$new_n1420 ;
  wire \$abc$9276$new_n1421 ;
  wire \$abc$9276$new_n1422 ;
  wire \$abc$9276$new_n1423 ;
  wire \$abc$9276$new_n1424 ;
  wire \$abc$9276$new_n1426 ;
  wire \$abc$9276$new_n1428 ;
  wire \$abc$9276$new_n1429 ;
  wire \$abc$9276$new_n1430 ;
  wire \$abc$9276$new_n1431 ;
  wire \$abc$9276$new_n1432 ;
  wire \$abc$9276$new_n1433 ;
  wire \$abc$9276$new_n1434 ;
  wire \$abc$9276$new_n1435 ;
  wire \$abc$9276$new_n1436 ;
  wire \$abc$9276$new_n1437 ;
  wire \$abc$9276$new_n1438 ;
  wire \$abc$9276$new_n1439 ;
  wire \$abc$9276$new_n1440 ;
  wire \$abc$9276$new_n1441 ;
  wire \$abc$9276$new_n1442 ;
  wire \$abc$9276$new_n1443 ;
  wire \$abc$9276$new_n1444 ;
  wire \$abc$9276$new_n1445 ;
  wire \$abc$9276$new_n1446 ;
  wire \$abc$9276$new_n1447 ;
  wire \$abc$9276$new_n1448 ;
  wire \$abc$9276$new_n1449 ;
  wire \$abc$9276$new_n1450 ;
  wire \$abc$9276$new_n1451 ;
  wire \$abc$9276$new_n1452 ;
  wire \$abc$9276$new_n1453 ;
  wire \$abc$9276$new_n1454 ;
  wire \$abc$9276$new_n1455 ;
  wire \$abc$9276$new_n1456 ;
  wire \$abc$9276$new_n1457 ;
  wire \$abc$9276$new_n1458 ;
  wire \$abc$9276$new_n1459 ;
  wire \$abc$9276$new_n1460 ;
  wire \$abc$9276$new_n1461 ;
  wire \$abc$9276$new_n1462 ;
  wire \$abc$9276$new_n1463 ;
  wire \$abc$9276$new_n1464 ;
  wire \$abc$9276$new_n1465 ;
  wire \$abc$9276$new_n1466 ;
  wire \$abc$9276$new_n1467 ;
  wire \$abc$9276$new_n1468 ;
  wire \$abc$9276$new_n1469 ;
  wire \$abc$9276$new_n1470 ;
  wire \$abc$9276$new_n1471 ;
  wire \$abc$9276$new_n1472 ;
  wire \$abc$9276$new_n1473 ;
  wire \$abc$9276$new_n1474 ;
  wire \$abc$9276$new_n1475 ;
  wire \$abc$9276$new_n1476 ;
  wire \$abc$9276$new_n1477 ;
  wire \$abc$9276$new_n1478 ;
  wire \$abc$9276$new_n1479 ;
  wire \$abc$9276$new_n1480 ;
  wire \$abc$9276$new_n1481 ;
  wire \$abc$9276$new_n1482 ;
  wire \$abc$9276$new_n1483 ;
  wire \$abc$9276$new_n1484 ;
  wire \$abc$9276$new_n1485 ;
  wire \$abc$9276$new_n1486 ;
  wire \$abc$9276$new_n1487 ;
  wire \$abc$9276$new_n1488 ;
  wire \$abc$9276$new_n1489 ;
  wire \$abc$9276$new_n1490 ;
  wire \$abc$9276$new_n1491 ;
  wire \$abc$9276$new_n1492 ;
  wire \$abc$9276$new_n1493 ;
  wire \$abc$9276$new_n1494 ;
  wire \$abc$9276$new_n1495 ;
  wire \$abc$9276$new_n1496 ;
  wire \$abc$9276$new_n1497 ;
  wire \$abc$9276$new_n1498 ;
  wire \$abc$9276$new_n1499 ;
  wire \$abc$9276$new_n1500 ;
  wire \$abc$9276$new_n1502 ;
  wire \$abc$9276$new_n1503 ;
  wire \$abc$9276$new_n1504 ;
  wire \$abc$9276$new_n1505 ;
  wire \$abc$9276$new_n1506 ;
  wire \$abc$9276$new_n1507 ;
  wire \$abc$9276$new_n1508 ;
  wire \$abc$9276$new_n1509 ;
  wire \$abc$9276$new_n1510 ;
  wire \$abc$9276$new_n1511 ;
  wire \$abc$9276$new_n1513 ;
  wire \$abc$9276$new_n1514 ;
  wire \$abc$9276$new_n1515 ;
  wire \$abc$9276$new_n1516 ;
  wire \$abc$9276$new_n1517 ;
  wire \$abc$9276$new_n1518 ;
  wire \$abc$9276$new_n1519 ;
  wire \$abc$9276$new_n1520 ;
  wire \$abc$9276$new_n1521 ;
  wire \$abc$9276$new_n1522 ;
  wire \$abc$9276$new_n1523 ;
  wire \$abc$9276$new_n1524 ;
  wire \$abc$9276$new_n1525 ;
  wire \$abc$9276$new_n1526 ;
  wire \$abc$9276$new_n1527 ;
  wire \$abc$9276$new_n1528 ;
  wire \$abc$9276$new_n1529 ;
  wire \$abc$9276$new_n1530 ;
  wire \$abc$9276$new_n1531 ;
  wire \$abc$9276$new_n1533 ;
  wire \$abc$9276$new_n1534 ;
  wire \$abc$9276$new_n1536 ;
  wire \$abc$9276$new_n1537 ;
  wire \$abc$9276$new_n1538 ;
  wire \$abc$9276$new_n1539 ;
  wire \$abc$9276$new_n1540 ;
  wire \$abc$9276$new_n1541 ;
  wire \$abc$9276$new_n1542 ;
  wire \$abc$9276$new_n1543 ;
  wire \$abc$9276$new_n1544 ;
  wire \$abc$9276$new_n1545 ;
  wire \$abc$9276$new_n1546 ;
  wire \$abc$9276$new_n1547 ;
  wire \$abc$9276$new_n1548 ;
  wire \$abc$9276$new_n1549 ;
  wire \$abc$9276$new_n1550 ;
  wire \$abc$9276$new_n1551 ;
  wire \$abc$9276$new_n1552 ;
  wire \$abc$9276$new_n1553 ;
  wire \$abc$9276$new_n1554 ;
  wire \$abc$9276$new_n1555 ;
  wire \$abc$9276$new_n1556 ;
  wire \$abc$9276$new_n1558 ;
  wire \$abc$9276$new_n1559 ;
  wire \$abc$9276$new_n1561 ;
  wire \$abc$9276$new_n1562 ;
  wire \$abc$9276$new_n1563 ;
  wire \$abc$9276$new_n1564 ;
  wire \$abc$9276$new_n1565 ;
  wire \$abc$9276$new_n1566 ;
  wire \$abc$9276$new_n1567 ;
  wire \$abc$9276$new_n1568 ;
  wire \$abc$9276$new_n1569 ;
  wire \$abc$9276$new_n1570 ;
  wire \$abc$9276$new_n1571 ;
  wire \$abc$9276$new_n1572 ;
  wire \$abc$9276$new_n1573 ;
  wire \$abc$9276$new_n1574 ;
  wire \$abc$9276$new_n1575 ;
  wire \$abc$9276$new_n1576 ;
  wire \$abc$9276$new_n1577 ;
  wire \$abc$9276$new_n1578 ;
  wire \$abc$9276$new_n1579 ;
  wire \$abc$9276$new_n1580 ;
  wire \$abc$9276$new_n1581 ;
  wire \$abc$9276$new_n1582 ;
  wire \$abc$9276$new_n1584 ;
  wire \$abc$9276$new_n1585 ;
  wire \$abc$9276$new_n1587 ;
  wire \$abc$9276$new_n1588 ;
  wire \$abc$9276$new_n1589 ;
  wire \$abc$9276$new_n1590 ;
  wire \$abc$9276$new_n1591 ;
  wire \$abc$9276$new_n1592 ;
  wire \$abc$9276$new_n1593 ;
  wire \$abc$9276$new_n1594 ;
  wire \$abc$9276$new_n1595 ;
  wire \$abc$9276$new_n1596 ;
  wire \$abc$9276$new_n1597 ;
  wire \$abc$9276$new_n1598 ;
  wire \$abc$9276$new_n1599 ;
  wire \$abc$9276$new_n1600 ;
  wire \$abc$9276$new_n1601 ;
  wire \$abc$9276$new_n1602 ;
  wire \$abc$9276$new_n1603 ;
  wire \$abc$9276$new_n1604 ;
  wire \$abc$9276$new_n1605 ;
  wire \$abc$9276$new_n1606 ;
  wire \$abc$9276$new_n1607 ;
  wire \$abc$9276$new_n1608 ;
  wire \$abc$9276$new_n1610 ;
  wire \$abc$9276$new_n1611 ;
  wire \$abc$9276$new_n1613 ;
  wire \$abc$9276$new_n1614 ;
  wire \$abc$9276$new_n1615 ;
  wire \$abc$9276$new_n1616 ;
  wire \$abc$9276$new_n1617 ;
  wire \$abc$9276$new_n1618 ;
  wire \$abc$9276$new_n1619 ;
  wire \$abc$9276$new_n1620 ;
  wire \$abc$9276$new_n1621 ;
  wire \$abc$9276$new_n1622 ;
  wire \$abc$9276$new_n1623 ;
  wire \$abc$9276$new_n1624 ;
  wire \$abc$9276$new_n1625 ;
  wire \$abc$9276$new_n1626 ;
  wire \$abc$9276$new_n1627 ;
  wire \$abc$9276$new_n1628 ;
  wire \$abc$9276$new_n1629 ;
  wire \$abc$9276$new_n1630 ;
  wire \$abc$9276$new_n1631 ;
  wire \$abc$9276$new_n1632 ;
  wire \$abc$9276$new_n1633 ;
  wire \$abc$9276$new_n1634 ;
  wire \$abc$9276$new_n1636 ;
  wire \$abc$9276$new_n1637 ;
  wire \$abc$9276$new_n1639 ;
  wire \$abc$9276$new_n1640 ;
  wire \$abc$9276$new_n1641 ;
  wire \$abc$9276$new_n1642 ;
  wire \$abc$9276$new_n1643 ;
  wire \$abc$9276$new_n1644 ;
  wire \$abc$9276$new_n1645 ;
  wire \$abc$9276$new_n1646 ;
  wire \$abc$9276$new_n1647 ;
  wire \$abc$9276$new_n1648 ;
  wire \$abc$9276$new_n1649 ;
  wire \$abc$9276$new_n1650 ;
  wire \$abc$9276$new_n1651 ;
  wire \$abc$9276$new_n1652 ;
  wire \$abc$9276$new_n1653 ;
  wire \$abc$9276$new_n1654 ;
  wire \$abc$9276$new_n1655 ;
  wire \$abc$9276$new_n1656 ;
  wire \$abc$9276$new_n1657 ;
  wire \$abc$9276$new_n1658 ;
  wire \$abc$9276$new_n1659 ;
  wire \$abc$9276$new_n1660 ;
  wire \$abc$9276$new_n1662 ;
  wire \$abc$9276$new_n1663 ;
  wire \$abc$9276$new_n1665 ;
  wire \$abc$9276$new_n1666 ;
  wire \$abc$9276$new_n1667 ;
  wire \$abc$9276$new_n1668 ;
  wire \$abc$9276$new_n1669 ;
  wire \$abc$9276$new_n1670 ;
  wire \$abc$9276$new_n1671 ;
  wire \$abc$9276$new_n1672 ;
  wire \$abc$9276$new_n1673 ;
  wire \$abc$9276$new_n1674 ;
  wire \$abc$9276$new_n1675 ;
  wire \$abc$9276$new_n1676 ;
  wire \$abc$9276$new_n1677 ;
  wire \$abc$9276$new_n1678 ;
  wire \$abc$9276$new_n1679 ;
  wire \$abc$9276$new_n1680 ;
  wire \$abc$9276$new_n1681 ;
  wire \$abc$9276$new_n1682 ;
  wire \$abc$9276$new_n1683 ;
  wire \$abc$9276$new_n1684 ;
  wire \$abc$9276$new_n1686 ;
  wire \$abc$9276$new_n1687 ;
  wire \$abc$9276$new_n1689 ;
  wire \$abc$9276$new_n1690 ;
  wire \$abc$9276$new_n1691 ;
  wire \$abc$9276$new_n1692 ;
  wire \$abc$9276$new_n1693 ;
  wire \$abc$9276$new_n1694 ;
  wire \$abc$9276$new_n1695 ;
  wire \$abc$9276$new_n1696 ;
  wire \$abc$9276$new_n1697 ;
  wire \$abc$9276$new_n1698 ;
  wire \$abc$9276$new_n1700 ;
  wire \$abc$9276$new_n1701 ;
  wire \$abc$9276$new_n1703 ;
  wire \$abc$9276$new_n1704 ;
  wire \$abc$9276$new_n1705 ;
  wire \$abc$9276$new_n1706 ;
  wire \$abc$9276$new_n1707 ;
  wire \$abc$9276$new_n1708 ;
  wire \$abc$9276$new_n1709 ;
  wire \$abc$9276$new_n1710 ;
  wire \$abc$9276$new_n1712 ;
  wire \$abc$9276$new_n1713 ;
  wire \$abc$9276$new_n1715 ;
  wire \$abc$9276$new_n1716 ;
  wire \$abc$9276$new_n1717 ;
  wire \$abc$9276$new_n1718 ;
  wire \$abc$9276$new_n1719 ;
  wire \$abc$9276$new_n1720 ;
  wire \$abc$9276$new_n1721 ;
  wire \$abc$9276$new_n1722 ;
  wire \$abc$9276$new_n1724 ;
  wire \$abc$9276$new_n1725 ;
  wire \$abc$9276$new_n1727 ;
  wire \$abc$9276$new_n1728 ;
  wire \$abc$9276$new_n1729 ;
  wire \$abc$9276$new_n1730 ;
  wire \$abc$9276$new_n1731 ;
  wire \$abc$9276$new_n1732 ;
  wire \$abc$9276$new_n1733 ;
  wire \$abc$9276$new_n1734 ;
  wire \$abc$9276$new_n1736 ;
  wire \$abc$9276$new_n1737 ;
  wire \$abc$9276$new_n1739 ;
  wire \$abc$9276$new_n1740 ;
  wire \$abc$9276$new_n1741 ;
  wire \$abc$9276$new_n1742 ;
  wire \$abc$9276$new_n1743 ;
  wire \$abc$9276$new_n1744 ;
  wire \$abc$9276$new_n1745 ;
  wire \$abc$9276$new_n1746 ;
  wire \$abc$9276$new_n1748 ;
  wire \$abc$9276$new_n1749 ;
  wire \$abc$9276$new_n1751 ;
  wire \$abc$9276$new_n1752 ;
  wire \$abc$9276$new_n1753 ;
  wire \$abc$9276$new_n1754 ;
  wire \$abc$9276$new_n1755 ;
  wire \$abc$9276$new_n1756 ;
  wire \$abc$9276$new_n1757 ;
  wire \$abc$9276$new_n1758 ;
  wire \$abc$9276$new_n1760 ;
  wire \$abc$9276$new_n1761 ;
  wire \$abc$9276$new_n1763 ;
  wire \$abc$9276$new_n1764 ;
  wire \$abc$9276$new_n1765 ;
  wire \$abc$9276$new_n1766 ;
  wire \$abc$9276$new_n1767 ;
  wire \$abc$9276$new_n1768 ;
  wire \$abc$9276$new_n1769 ;
  wire \$abc$9276$new_n1770 ;
  wire \$abc$9276$new_n1771 ;
  wire \$abc$9276$new_n1772 ;
  wire \$abc$9276$new_n1774 ;
  wire \$abc$9276$new_n1775 ;
  wire \$abc$9276$new_n1777 ;
  wire \$abc$9276$new_n1778 ;
  wire \$abc$9276$new_n1779 ;
  wire \$abc$9276$new_n1780 ;
  wire \$abc$9276$new_n1781 ;
  wire \$abc$9276$new_n1782 ;
  wire \$abc$9276$new_n1783 ;
  wire \$abc$9276$new_n1784 ;
  wire \$abc$9276$new_n1786 ;
  wire \$abc$9276$new_n1787 ;
  wire \$abc$9276$new_n1789 ;
  wire \$abc$9276$new_n1790 ;
  wire \$abc$9276$new_n1791 ;
  wire \$abc$9276$new_n1792 ;
  wire \$abc$9276$new_n1793 ;
  wire \$abc$9276$new_n1795 ;
  wire \$abc$9276$new_n1796 ;
  wire \$abc$9276$new_n1798 ;
  wire \$abc$9276$new_n1799 ;
  wire \$abc$9276$new_n1801 ;
  wire \$abc$9276$new_n1802 ;
  wire \$abc$9276$new_n1804 ;
  wire \$abc$9276$new_n1805 ;
  wire \$abc$9276$new_n1807 ;
  wire \$abc$9276$new_n1808 ;
  wire \$abc$9276$new_n1810 ;
  wire \$abc$9276$new_n1811 ;
  wire \$abc$9276$new_n1813 ;
  wire \$abc$9276$new_n1814 ;
  wire \$abc$9276$new_n1816 ;
  wire \$abc$9276$new_n1817 ;
  wire \$abc$9276$new_n1818 ;
  wire \$abc$9276$new_n1819 ;
  wire \$abc$9276$new_n1820 ;
  wire \$abc$9276$new_n1821 ;
  wire \$abc$9276$new_n1822 ;
  wire \$abc$9276$new_n1823 ;
  wire \$abc$9276$new_n1824 ;
  wire \$abc$9276$new_n1825 ;
  wire \$abc$9276$new_n1826 ;
  wire \$abc$9276$new_n1827 ;
  wire \$abc$9276$new_n1828 ;
  wire \$abc$9276$new_n1829 ;
  wire \$abc$9276$new_n1830 ;
  wire \$abc$9276$new_n1831 ;
  wire \$abc$9276$new_n1832 ;
  wire \$abc$9276$new_n1833 ;
  wire \$abc$9276$new_n1834 ;
  wire \$abc$9276$new_n1835 ;
  wire \$abc$9276$new_n1836 ;
  wire \$abc$9276$new_n1837 ;
  wire \$abc$9276$new_n1838 ;
  wire \$abc$9276$new_n1839 ;
  wire \$abc$9276$new_n1840 ;
  wire \$abc$9276$new_n1841 ;
  wire \$abc$9276$new_n1842 ;
  wire \$abc$9276$new_n1843 ;
  wire \$abc$9276$new_n1844 ;
  wire \$abc$9276$new_n1845 ;
  wire \$abc$9276$new_n1846 ;
  wire \$abc$9276$new_n1847 ;
  wire \$abc$9276$new_n1848 ;
  wire \$abc$9276$new_n1849 ;
  wire \$abc$9276$new_n1850 ;
  wire \$abc$9276$new_n1851 ;
  wire \$abc$9276$new_n1852 ;
  wire \$abc$9276$new_n1853 ;
  wire \$abc$9276$new_n1854 ;
  wire \$abc$9276$new_n1855 ;
  wire \$abc$9276$new_n1856 ;
  wire \$abc$9276$new_n1857 ;
  wire \$abc$9276$new_n1858 ;
  wire \$abc$9276$new_n1859 ;
  wire \$abc$9276$new_n1860 ;
  wire \$abc$9276$new_n1861 ;
  wire \$abc$9276$new_n1862 ;
  wire \$abc$9276$new_n1863 ;
  wire \$abc$9276$new_n1864 ;
  wire \$abc$9276$new_n1865 ;
  wire \$abc$9276$new_n1866 ;
  wire \$abc$9276$new_n1867 ;
  wire \$abc$9276$new_n1868 ;
  wire \$abc$9276$new_n1869 ;
  wire \$abc$9276$new_n1870 ;
  wire \$abc$9276$new_n1871 ;
  wire \$abc$9276$new_n1872 ;
  wire \$abc$9276$new_n1873 ;
  wire \$abc$9276$new_n1874 ;
  wire \$abc$9276$new_n1875 ;
  wire \$abc$9276$new_n1876 ;
  wire \$abc$9276$new_n1877 ;
  wire \$abc$9276$new_n1878 ;
  wire \$abc$9276$new_n1879 ;
  wire \$abc$9276$new_n1880 ;
  wire \$abc$9276$new_n1881 ;
  wire \$abc$9276$new_n1882 ;
  wire \$abc$9276$new_n1883 ;
  wire \$abc$9276$new_n1884 ;
  wire \$abc$9276$new_n1885 ;
  wire \$abc$9276$new_n1886 ;
  wire \$abc$9276$new_n1887 ;
  wire \$abc$9276$new_n1888 ;
  wire \$abc$9276$new_n1889 ;
  wire \$abc$9276$new_n1890 ;
  wire \$abc$9276$new_n1891 ;
  wire \$abc$9276$new_n1892 ;
  wire \$abc$9276$new_n1893 ;
  wire \$abc$9276$new_n1894 ;
  wire \$abc$9276$new_n1895 ;
  wire \$abc$9276$new_n1896 ;
  wire \$abc$9276$new_n1897 ;
  wire \$abc$9276$new_n1898 ;
  wire \$abc$9276$new_n1899 ;
  wire \$abc$9276$new_n1900 ;
  wire \$abc$9276$new_n1901 ;
  wire \$abc$9276$new_n1902 ;
  wire \$abc$9276$new_n1903 ;
  wire \$abc$9276$new_n1904 ;
  wire \$abc$9276$new_n1905 ;
  wire \$abc$9276$new_n1906 ;
  wire \$abc$9276$new_n1907 ;
  wire \$abc$9276$new_n1908 ;
  wire \$abc$9276$new_n1909 ;
  wire \$abc$9276$new_n1910 ;
  wire \$abc$9276$new_n1911 ;
  wire \$abc$9276$new_n1912 ;
  wire \$abc$9276$new_n1913 ;
  wire \$abc$9276$new_n1914 ;
  wire \$abc$9276$new_n1915 ;
  wire \$abc$9276$new_n1916 ;
  wire \$abc$9276$new_n1917 ;
  wire \$abc$9276$new_n1918 ;
  wire \$abc$9276$new_n1919 ;
  wire \$abc$9276$new_n1920 ;
  wire \$abc$9276$new_n1921 ;
  wire \$abc$9276$new_n1922 ;
  wire \$abc$9276$new_n1923 ;
  wire \$abc$9276$new_n1924 ;
  wire \$abc$9276$new_n1925 ;
  wire \$abc$9276$new_n1926 ;
  wire \$abc$9276$new_n1927 ;
  wire \$abc$9276$new_n1928 ;
  wire \$abc$9276$new_n1929 ;
  wire \$abc$9276$new_n1930 ;
  wire \$abc$9276$new_n1931 ;
  wire \$abc$9276$new_n1932 ;
  wire \$abc$9276$new_n1933 ;
  wire \$abc$9276$new_n1934 ;
  wire \$abc$9276$new_n1935 ;
  wire \$abc$9276$new_n1936 ;
  wire \$abc$9276$new_n1937 ;
  wire \$abc$9276$new_n1938 ;
  wire \$abc$9276$new_n1939 ;
  wire \$abc$9276$new_n1940 ;
  wire \$abc$9276$new_n1941 ;
  wire \$abc$9276$new_n1942 ;
  wire \$abc$9276$new_n1943 ;
  wire \$abc$9276$new_n1945 ;
  wire \$abc$9276$new_n1946 ;
  wire \$abc$9276$new_n1947 ;
  wire \$abc$9276$new_n1948 ;
  wire \$abc$9276$new_n1949 ;
  wire \$abc$9276$new_n1950 ;
  wire \$abc$9276$new_n1951 ;
  wire \$abc$9276$new_n1952 ;
  wire \$abc$9276$new_n1953 ;
  wire \$abc$9276$new_n1954 ;
  wire \$abc$9276$new_n1955 ;
  wire \$abc$9276$new_n1956 ;
  wire \$abc$9276$new_n1957 ;
  wire \$abc$9276$new_n1958 ;
  wire \$abc$9276$new_n1959 ;
  wire \$abc$9276$new_n1960 ;
  wire \$abc$9276$new_n1961 ;
  wire \$abc$9276$new_n1962 ;
  wire \$abc$9276$new_n1963 ;
  wire \$abc$9276$new_n1964 ;
  wire \$abc$9276$new_n1965 ;
  wire \$abc$9276$new_n1966 ;
  wire \$abc$9276$new_n1967 ;
  wire \$abc$9276$new_n1968 ;
  wire \$abc$9276$new_n1969 ;
  wire \$abc$9276$new_n1970 ;
  wire \$abc$9276$new_n1971 ;
  wire \$abc$9276$new_n1972 ;
  wire \$abc$9276$new_n1973 ;
  wire \$abc$9276$new_n1974 ;
  wire \$abc$9276$new_n1975 ;
  wire \$abc$9276$new_n1976 ;
  wire \$abc$9276$new_n1977 ;
  wire \$abc$9276$new_n1978 ;
  wire \$abc$9276$new_n1979 ;
  wire \$abc$9276$new_n1980 ;
  wire \$abc$9276$new_n1981 ;
  wire \$abc$9276$new_n1982 ;
  wire \$abc$9276$new_n1983 ;
  wire \$abc$9276$new_n1984 ;
  wire \$abc$9276$new_n1985 ;
  wire \$abc$9276$new_n1986 ;
  wire \$abc$9276$new_n1987 ;
  wire \$abc$9276$new_n1988 ;
  wire \$abc$9276$new_n1989 ;
  wire \$abc$9276$new_n1990 ;
  wire \$abc$9276$new_n1991 ;
  wire \$abc$9276$new_n1992 ;
  wire \$abc$9276$new_n1993 ;
  wire \$abc$9276$new_n1994 ;
  wire \$abc$9276$new_n1995 ;
  wire \$abc$9276$new_n1996 ;
  wire \$abc$9276$new_n1997 ;
  wire \$abc$9276$new_n1998 ;
  wire \$abc$9276$new_n2000 ;
  wire \$abc$9276$new_n2001 ;
  wire \$abc$9276$new_n2002 ;
  wire \$abc$9276$new_n2003 ;
  wire \$abc$9276$new_n2004 ;
  wire \$abc$9276$new_n2005 ;
  wire \$abc$9276$new_n2006 ;
  wire \$abc$9276$new_n2007 ;
  wire \$abc$9276$new_n2008 ;
  wire \$abc$9276$new_n2009 ;
  wire \$abc$9276$new_n2010 ;
  wire \$abc$9276$new_n2011 ;
  wire \$abc$9276$new_n2012 ;
  wire \$abc$9276$new_n2013 ;
  wire \$abc$9276$new_n2014 ;
  wire \$abc$9276$new_n2015 ;
  wire \$abc$9276$new_n2016 ;
  wire \$abc$9276$new_n2017 ;
  wire \$abc$9276$new_n2018 ;
  wire \$abc$9276$new_n2019 ;
  wire \$abc$9276$new_n2020 ;
  wire \$abc$9276$new_n2021 ;
  wire \$abc$9276$new_n2022 ;
  wire \$abc$9276$new_n2024 ;
  wire \$abc$9276$new_n2025 ;
  wire \$abc$9276$new_n2026 ;
  wire \$abc$9276$new_n2027 ;
  wire \$abc$9276$new_n2028 ;
  wire \$abc$9276$new_n2029 ;
  wire \$abc$9276$new_n2030 ;
  wire \$abc$9276$new_n2031 ;
  wire \$abc$9276$new_n2032 ;
  wire \$abc$9276$new_n2033 ;
  wire \$abc$9276$new_n2034 ;
  wire \$abc$9276$new_n2035 ;
  wire \$abc$9276$new_n2036 ;
  wire \$abc$9276$new_n2037 ;
  wire \$abc$9276$new_n2038 ;
  wire \$abc$9276$new_n2039 ;
  wire \$abc$9276$new_n2040 ;
  wire \$abc$9276$new_n2041 ;
  wire \$abc$9276$new_n2042 ;
  wire \$abc$9276$new_n2043 ;
  wire \$abc$9276$new_n2044 ;
  wire \$abc$9276$new_n2045 ;
  wire \$abc$9276$new_n2046 ;
  wire \$abc$9276$new_n2047 ;
  wire \$abc$9276$new_n2048 ;
  wire \$abc$9276$new_n2049 ;
  wire \$abc$9276$new_n2051 ;
  wire \$abc$9276$new_n2052 ;
  wire \$abc$9276$new_n2053 ;
  wire \$abc$9276$new_n2054 ;
  wire \$abc$9276$new_n2055 ;
  wire \$abc$9276$new_n2056 ;
  wire \$abc$9276$new_n2057 ;
  wire \$abc$9276$new_n2058 ;
  wire \$abc$9276$new_n2059 ;
  wire \$abc$9276$new_n2060 ;
  wire \$abc$9276$new_n2061 ;
  wire \$abc$9276$new_n2062 ;
  wire \$abc$9276$new_n2063 ;
  wire \$abc$9276$new_n2064 ;
  wire \$abc$9276$new_n2065 ;
  wire \$abc$9276$new_n2066 ;
  wire \$abc$9276$new_n2067 ;
  wire \$abc$9276$new_n2068 ;
  wire \$abc$9276$new_n2070 ;
  wire \$abc$9276$new_n2071 ;
  wire \$abc$9276$new_n2072 ;
  wire \$abc$9276$new_n2073 ;
  wire \$abc$9276$new_n2074 ;
  wire \$abc$9276$new_n2075 ;
  wire \$abc$9276$new_n2076 ;
  wire \$abc$9276$new_n2077 ;
  wire \$abc$9276$new_n2078 ;
  wire \$abc$9276$new_n2079 ;
  wire \$abc$9276$new_n2080 ;
  wire \$abc$9276$new_n2081 ;
  wire \$abc$9276$new_n2082 ;
  wire \$abc$9276$new_n2084 ;
  wire \$abc$9276$new_n2085 ;
  wire \$abc$9276$new_n2086 ;
  wire \$abc$9276$new_n2087 ;
  wire \$abc$9276$new_n2088 ;
  wire \$abc$9276$new_n2089 ;
  wire \$abc$9276$new_n2090 ;
  wire \$abc$9276$new_n2091 ;
  wire \$abc$9276$new_n2092 ;
  wire \$abc$9276$new_n2093 ;
  wire \$abc$9276$new_n2094 ;
  wire \$abc$9276$new_n2095 ;
  wire \$abc$9276$new_n2096 ;
  wire \$abc$9276$new_n2097 ;
  wire \$abc$9276$new_n2098 ;
  wire \$abc$9276$new_n2100 ;
  wire \$abc$9276$new_n2101 ;
  wire \$abc$9276$new_n2102 ;
  wire \$abc$9276$new_n2103 ;
  wire \$abc$9276$new_n2104 ;
  wire \$abc$9276$new_n2105 ;
  wire \$abc$9276$new_n2106 ;
  wire \$abc$9276$new_n2107 ;
  wire \$abc$9276$new_n2109 ;
  wire \$abc$9276$new_n2110 ;
  wire \$abc$9276$new_n2111 ;
  wire \$abc$9276$new_n2112 ;
  wire \$abc$9276$new_n2113 ;
  wire \$abc$9276$new_n2114 ;
  wire \$abc$9276$new_n2115 ;
  wire \$abc$9276$new_n2116 ;
  wire \$abc$9276$new_n2117 ;
  wire \$abc$9276$new_n2118 ;
  wire \$abc$9276$new_n2119 ;
  wire \$abc$9276$new_n2120 ;
  wire \$abc$9276$new_n2121 ;
  wire \$abc$9276$new_n2122 ;
  wire \$abc$9276$new_n2123 ;
  wire \$abc$9276$new_n2124 ;
  wire \$abc$9276$new_n2125 ;
  wire \$abc$9276$new_n2127 ;
  wire \$abc$9276$new_n2128 ;
  wire \$abc$9276$new_n2129 ;
  wire \$abc$9276$new_n2130 ;
  wire \$abc$9276$new_n2131 ;
  wire \$abc$9276$new_n2133 ;
  wire \$abc$9276$new_n2134 ;
  wire \$abc$9276$new_n2135 ;
  wire \$abc$9276$new_n2136 ;
  wire \$abc$9276$new_n2137 ;
  wire \$abc$9276$new_n2138 ;
  wire \$abc$9276$new_n2139 ;
  wire \$abc$9276$new_n2140 ;
  wire \$abc$9276$new_n2141 ;
  wire \$abc$9276$new_n2142 ;
  wire \$abc$9276$new_n2143 ;
  wire \$abc$9276$new_n2144 ;
  wire \$abc$9276$new_n2145 ;
  wire \$abc$9276$new_n2147 ;
  wire \$abc$9276$new_n2148 ;
  wire \$abc$9276$new_n2149 ;
  wire \$abc$9276$new_n2150 ;
  wire \$abc$9276$new_n2151 ;
  wire \$abc$9276$new_n2152 ;
  wire \$abc$9276$new_n2153 ;
  wire \$abc$9276$new_n2154 ;
  wire \$abc$9276$new_n2155 ;
  wire \$abc$9276$new_n2156 ;
  wire \$abc$9276$new_n2157 ;
  wire \$abc$9276$new_n2158 ;
  wire \$abc$9276$new_n2160 ;
  wire \$abc$9276$new_n2161 ;
  wire \$abc$9276$new_n2162 ;
  wire \$abc$9276$new_n2163 ;
  wire \$abc$9276$new_n2164 ;
  wire \$abc$9276$new_n2165 ;
  wire \$abc$9276$new_n2166 ;
  wire \$abc$9276$new_n2167 ;
  wire \$abc$9276$new_n2168 ;
  wire \$abc$9276$new_n2170 ;
  wire \$abc$9276$new_n2171 ;
  wire \$abc$9276$new_n2172 ;
  wire \$abc$9276$new_n2173 ;
  wire \$abc$9276$new_n2174 ;
  wire \$abc$9276$new_n2175 ;
  wire \$abc$9276$new_n2177 ;
  wire \$abc$9276$new_n2178 ;
  wire \$abc$9276$new_n2179 ;
  wire \$abc$9276$new_n2180 ;
  wire \$abc$9276$new_n2181 ;
  wire \$abc$9276$new_n2182 ;
  wire \$abc$9276$new_n2183 ;
  wire \$abc$9276$new_n2184 ;
  wire \$abc$9276$new_n2185 ;
  wire \$abc$9276$new_n2186 ;
  wire \$abc$9276$new_n2187 ;
  wire \$abc$9276$new_n2188 ;
  wire \$abc$9276$new_n2189 ;
  wire \$abc$9276$new_n2190 ;
  wire \$abc$9276$new_n2191 ;
  wire \$abc$9276$new_n2192 ;
  wire \$abc$9276$new_n2193 ;
  wire \$abc$9276$new_n2194 ;
  wire \$abc$9276$new_n2195 ;
  wire \$abc$9276$new_n2196 ;
  wire \$abc$9276$new_n2197 ;
  wire \$abc$9276$new_n2198 ;
  wire \$abc$9276$new_n2199 ;
  wire \$abc$9276$new_n2200 ;
  wire \$abc$9276$new_n2201 ;
  wire \$abc$9276$new_n2202 ;
  wire \$abc$9276$new_n2203 ;
  wire \$abc$9276$new_n2204 ;
  wire \$abc$9276$new_n2205 ;
  wire \$abc$9276$new_n2206 ;
  wire \$abc$9276$new_n2207 ;
  wire \$abc$9276$new_n2208 ;
  wire \$abc$9276$new_n2209 ;
  wire \$abc$9276$new_n2210 ;
  wire \$abc$9276$new_n2211 ;
  wire \$abc$9276$new_n2212 ;
  wire \$abc$9276$new_n2213 ;
  wire \$abc$9276$new_n2214 ;
  wire \$abc$9276$new_n2215 ;
  wire \$abc$9276$new_n2216 ;
  wire \$abc$9276$new_n2217 ;
  wire \$abc$9276$new_n2218 ;
  wire \$abc$9276$new_n2219 ;
  wire \$abc$9276$new_n2220 ;
  wire \$abc$9276$new_n2221 ;
  wire \$abc$9276$new_n2222 ;
  wire \$abc$9276$new_n2223 ;
  wire \$abc$9276$new_n2224 ;
  wire \$abc$9276$new_n2225 ;
  wire \$abc$9276$new_n2226 ;
  wire \$abc$9276$new_n2227 ;
  wire \$abc$9276$new_n2228 ;
  wire \$abc$9276$new_n2229 ;
  wire \$abc$9276$new_n2230 ;
  wire \$abc$9276$new_n2231 ;
  wire \$abc$9276$new_n2232 ;
  wire \$abc$9276$new_n2233 ;
  wire \$abc$9276$new_n2234 ;
  wire \$abc$9276$new_n2235 ;
  wire \$abc$9276$new_n2236 ;
  wire \$abc$9276$new_n2237 ;
  wire \$abc$9276$new_n2238 ;
  wire \$abc$9276$new_n2239 ;
  wire \$abc$9276$new_n2240 ;
  wire \$abc$9276$new_n2241 ;
  wire \$abc$9276$new_n2242 ;
  wire \$abc$9276$new_n2243 ;
  wire \$abc$9276$new_n2244 ;
  wire \$abc$9276$new_n2245 ;
  wire \$abc$9276$new_n2246 ;
  wire \$abc$9276$new_n2247 ;
  wire \$abc$9276$new_n2248 ;
  wire \$abc$9276$new_n2249 ;
  wire \$abc$9276$new_n2250 ;
  wire \$abc$9276$new_n2251 ;
  wire \$abc$9276$new_n2252 ;
  wire \$abc$9276$new_n2253 ;
  wire \$abc$9276$new_n2254 ;
  wire \$abc$9276$new_n2255 ;
  wire \$abc$9276$new_n2256 ;
  wire \$abc$9276$new_n2257 ;
  wire \$abc$9276$new_n2258 ;
  wire \$abc$9276$new_n2259 ;
  wire \$abc$9276$new_n2260 ;
  wire \$abc$9276$new_n2261 ;
  wire \$abc$9276$new_n2262 ;
  wire \$abc$9276$new_n2263 ;
  wire \$abc$9276$new_n2264 ;
  wire \$abc$9276$new_n2265 ;
  wire \$abc$9276$new_n2266 ;
  wire \$abc$9276$new_n2267 ;
  wire \$abc$9276$new_n2268 ;
  wire \$abc$9276$new_n2269 ;
  wire \$abc$9276$new_n2270 ;
  wire \$abc$9276$new_n2271 ;
  wire \$abc$9276$new_n2272 ;
  wire \$abc$9276$new_n2273 ;
  wire \$abc$9276$new_n2274 ;
  wire \$abc$9276$new_n2275 ;
  wire \$abc$9276$new_n2276 ;
  wire \$abc$9276$new_n2277 ;
  wire \$abc$9276$new_n2278 ;
  wire \$abc$9276$new_n2279 ;
  wire \$abc$9276$new_n2280 ;
  wire \$abc$9276$new_n2281 ;
  wire \$abc$9276$new_n2282 ;
  wire \$abc$9276$new_n2283 ;
  wire \$abc$9276$new_n2284 ;
  wire \$abc$9276$new_n2285 ;
  wire \$abc$9276$new_n2286 ;
  wire \$abc$9276$new_n2287 ;
  wire \$abc$9276$new_n2288 ;
  wire \$abc$9276$new_n2289 ;
  wire \$abc$9276$new_n2290 ;
  wire \$abc$9276$new_n2291 ;
  wire \$abc$9276$new_n2292 ;
  wire \$abc$9276$new_n2293 ;
  wire \$abc$9276$new_n2294 ;
  wire \$abc$9276$new_n2295 ;
  wire \$abc$9276$new_n2296 ;
  wire \$abc$9276$new_n2297 ;
  wire \$abc$9276$new_n2298 ;
  wire \$abc$9276$new_n2299 ;
  wire \$abc$9276$new_n2300 ;
  wire \$abc$9276$new_n2301 ;
  wire \$abc$9276$new_n2302 ;
  wire \$abc$9276$new_n2303 ;
  wire \$abc$9276$new_n2304 ;
  wire \$abc$9276$new_n2305 ;
  wire \$abc$9276$new_n2307 ;
  wire \$abc$9276$new_n2308 ;
  wire \$abc$9276$new_n2309 ;
  wire \$abc$9276$new_n2310 ;
  wire \$abc$9276$new_n2311 ;
  wire \$abc$9276$new_n2312 ;
  wire \$abc$9276$new_n2313 ;
  wire \$abc$9276$new_n2314 ;
  wire \$abc$9276$new_n2315 ;
  wire \$abc$9276$new_n2316 ;
  wire \$abc$9276$new_n2317 ;
  wire \$abc$9276$new_n2318 ;
  wire \$abc$9276$new_n2319 ;
  wire \$abc$9276$new_n2320 ;
  wire \$abc$9276$new_n2321 ;
  wire \$abc$9276$new_n2322 ;
  wire \$abc$9276$new_n2323 ;
  wire \$abc$9276$new_n2324 ;
  wire \$abc$9276$new_n2325 ;
  wire \$abc$9276$new_n2326 ;
  wire \$abc$9276$new_n2327 ;
  wire \$abc$9276$new_n2328 ;
  wire \$abc$9276$new_n2329 ;
  wire \$abc$9276$new_n2330 ;
  wire \$abc$9276$new_n2331 ;
  wire \$abc$9276$new_n2332 ;
  wire \$abc$9276$new_n2333 ;
  wire \$abc$9276$new_n2334 ;
  wire \$abc$9276$new_n2335 ;
  wire \$abc$9276$new_n2336 ;
  wire \$abc$9276$new_n2337 ;
  wire \$abc$9276$new_n2338 ;
  wire \$abc$9276$new_n2339 ;
  wire \$abc$9276$new_n2340 ;
  wire \$abc$9276$new_n2341 ;
  wire \$abc$9276$new_n2342 ;
  wire \$abc$9276$new_n2343 ;
  wire \$abc$9276$new_n2344 ;
  wire \$abc$9276$new_n2345 ;
  wire \$abc$9276$new_n2346 ;
  wire \$abc$9276$new_n2347 ;
  wire \$abc$9276$new_n2348 ;
  wire \$abc$9276$new_n2349 ;
  wire \$abc$9276$new_n2350 ;
  wire \$abc$9276$new_n2351 ;
  wire \$abc$9276$new_n2352 ;
  wire \$abc$9276$new_n2353 ;
  wire \$abc$9276$new_n2354 ;
  wire \$abc$9276$new_n2355 ;
  wire \$abc$9276$new_n2356 ;
  wire \$abc$9276$new_n2357 ;
  wire \$abc$9276$new_n2358 ;
  wire \$abc$9276$new_n2359 ;
  wire \$abc$9276$new_n2360 ;
  wire \$abc$9276$new_n2361 ;
  wire \$abc$9276$new_n2362 ;
  wire \$abc$9276$new_n2363 ;
  wire \$abc$9276$new_n2364 ;
  wire \$abc$9276$new_n2365 ;
  wire \$abc$9276$new_n2366 ;
  wire \$abc$9276$new_n2367 ;
  wire \$abc$9276$new_n2368 ;
  wire \$abc$9276$new_n2369 ;
  wire \$abc$9276$new_n2370 ;
  wire \$abc$9276$new_n2371 ;
  wire \$abc$9276$new_n2372 ;
  wire \$abc$9276$new_n2373 ;
  wire \$abc$9276$new_n2374 ;
  wire \$abc$9276$new_n2375 ;
  wire \$abc$9276$new_n2376 ;
  wire \$abc$9276$new_n2377 ;
  wire \$abc$9276$new_n2378 ;
  wire \$abc$9276$new_n2379 ;
  wire \$abc$9276$new_n2380 ;
  wire \$abc$9276$new_n2381 ;
  wire \$abc$9276$new_n2382 ;
  wire \$abc$9276$new_n2383 ;
  wire \$abc$9276$new_n2384 ;
  wire \$abc$9276$new_n2385 ;
  wire \$abc$9276$new_n2386 ;
  wire \$abc$9276$new_n2387 ;
  wire \$abc$9276$new_n2388 ;
  wire \$abc$9276$new_n2389 ;
  wire \$abc$9276$new_n2390 ;
  wire \$abc$9276$new_n2391 ;
  wire \$abc$9276$new_n2392 ;
  wire \$abc$9276$new_n2393 ;
  wire \$abc$9276$new_n2394 ;
  wire \$abc$9276$new_n2395 ;
  wire \$abc$9276$new_n2396 ;
  wire \$abc$9276$new_n2397 ;
  wire \$abc$9276$new_n2398 ;
  wire \$abc$9276$new_n2399 ;
  wire \$abc$9276$new_n2400 ;
  wire \$abc$9276$new_n2401 ;
  wire \$abc$9276$new_n2402 ;
  wire \$abc$9276$new_n2403 ;
  wire \$abc$9276$new_n2404 ;
  wire \$abc$9276$new_n2405 ;
  wire \$abc$9276$new_n2406 ;
  wire \$abc$9276$new_n2407 ;
  wire \$abc$9276$new_n2408 ;
  wire \$abc$9276$new_n2409 ;
  wire \$abc$9276$new_n2410 ;
  wire \$abc$9276$new_n2411 ;
  wire \$abc$9276$new_n2412 ;
  wire \$abc$9276$new_n2413 ;
  wire \$abc$9276$new_n2414 ;
  wire \$abc$9276$new_n2415 ;
  wire \$abc$9276$new_n2416 ;
  wire \$abc$9276$new_n2417 ;
  wire \$abc$9276$new_n2418 ;
  wire \$abc$9276$new_n2419 ;
  wire \$abc$9276$new_n2420 ;
  wire \$abc$9276$new_n2421 ;
  wire \$abc$9276$new_n2422 ;
  wire \$abc$9276$new_n2423 ;
  wire \$abc$9276$new_n2424 ;
  wire \$abc$9276$new_n2425 ;
  wire \$abc$9276$new_n2426 ;
  wire \$abc$9276$new_n2427 ;
  wire \$abc$9276$new_n2428 ;
  wire \$abc$9276$new_n2429 ;
  wire \$abc$9276$new_n2430 ;
  wire \$abc$9276$new_n2431 ;
  wire \$abc$9276$new_n2432 ;
  wire \$abc$9276$new_n2433 ;
  wire \$abc$9276$new_n2434 ;
  wire \$abc$9276$new_n2435 ;
  wire \$abc$9276$new_n2436 ;
  wire \$abc$9276$new_n2437 ;
  wire \$abc$9276$new_n2438 ;
  wire \$abc$9276$new_n2439 ;
  wire \$abc$9276$new_n2440 ;
  wire \$abc$9276$new_n2441 ;
  wire \$abc$9276$new_n2442 ;
  wire \$abc$9276$new_n2443 ;
  wire \$abc$9276$new_n2444 ;
  wire \$abc$9276$new_n2445 ;
  wire \$abc$9276$new_n2446 ;
  wire \$abc$9276$new_n2447 ;
  wire \$abc$9276$new_n2448 ;
  wire \$abc$9276$new_n2449 ;
  wire \$abc$9276$new_n2450 ;
  wire \$abc$9276$new_n2451 ;
  wire \$abc$9276$new_n2452 ;
  wire \$abc$9276$new_n2453 ;
  wire \$abc$9276$new_n2454 ;
  wire \$abc$9276$new_n2455 ;
  wire \$abc$9276$new_n2456 ;
  wire \$abc$9276$new_n2457 ;
  wire \$abc$9276$new_n2458 ;
  wire \$abc$9276$new_n2459 ;
  wire \$abc$9276$new_n2460 ;
  wire \$abc$9276$new_n2461 ;
  wire \$abc$9276$new_n2462 ;
  wire \$abc$9276$new_n2463 ;
  wire \$abc$9276$new_n2464 ;
  wire \$abc$9276$new_n2465 ;
  wire \$abc$9276$new_n2466 ;
  wire \$abc$9276$new_n2467 ;
  wire \$abc$9276$new_n2468 ;
  wire \$abc$9276$new_n2469 ;
  wire \$abc$9276$new_n2470 ;
  wire \$abc$9276$new_n2471 ;
  wire \$abc$9276$new_n2472 ;
  wire \$abc$9276$new_n2473 ;
  wire \$abc$9276$new_n2474 ;
  wire \$abc$9276$new_n2475 ;
  wire \$abc$9276$new_n2476 ;
  wire \$abc$9276$new_n2477 ;
  wire \$abc$9276$new_n2478 ;
  wire \$abc$9276$new_n2479 ;
  wire \$abc$9276$new_n2480 ;
  wire \$abc$9276$new_n2481 ;
  wire \$abc$9276$new_n2482 ;
  wire \$abc$9276$new_n2483 ;
  wire \$abc$9276$new_n2484 ;
  wire \$abc$9276$new_n2485 ;
  wire \$abc$9276$new_n2486 ;
  wire \$abc$9276$new_n2487 ;
  wire \$abc$9276$new_n2488 ;
  wire \$abc$9276$new_n2489 ;
  wire \$abc$9276$new_n2490 ;
  wire \$abc$9276$new_n2491 ;
  wire \$abc$9276$new_n2492 ;
  wire \$abc$9276$new_n2493 ;
  wire \$abc$9276$new_n2494 ;
  wire \$abc$9276$new_n2495 ;
  wire \$abc$9276$new_n2496 ;
  wire \$abc$9276$new_n2497 ;
  wire \$abc$9276$new_n2498 ;
  wire \$abc$9276$new_n2499 ;
  wire \$abc$9276$new_n2500 ;
  wire \$abc$9276$new_n2501 ;
  wire \$abc$9276$new_n2502 ;
  wire \$abc$9276$new_n2503 ;
  wire \$abc$9276$new_n2504 ;
  wire \$abc$9276$new_n2505 ;
  wire \$abc$9276$new_n2506 ;
  wire \$abc$9276$new_n2507 ;
  wire \$abc$9276$new_n2508 ;
  wire \$abc$9276$new_n2509 ;
  wire \$abc$9276$new_n2510 ;
  wire \$abc$9276$new_n2511 ;
  wire \$abc$9276$new_n2512 ;
  wire \$abc$9276$new_n2513 ;
  wire \$abc$9276$new_n2514 ;
  wire \$abc$9276$new_n2515 ;
  wire \$abc$9276$new_n2516 ;
  wire \$abc$9276$new_n2517 ;
  wire \$abc$9276$new_n2518 ;
  wire \$abc$9276$new_n2519 ;
  wire \$abc$9276$new_n2520 ;
  wire \$abc$9276$new_n2521 ;
  wire \$abc$9276$new_n2522 ;
  wire \$abc$9276$new_n2523 ;
  wire \$abc$9276$new_n2524 ;
  wire \$abc$9276$new_n2525 ;
  wire \$abc$9276$new_n2526 ;
  wire \$abc$9276$new_n2527 ;
  wire \$abc$9276$new_n2528 ;
  wire \$abc$9276$new_n2529 ;
  wire \$abc$9276$new_n2530 ;
  wire \$abc$9276$new_n2531 ;
  wire \$abc$9276$new_n2532 ;
  wire \$abc$9276$new_n2533 ;
  wire \$abc$9276$new_n2534 ;
  wire \$abc$9276$new_n2535 ;
  wire \$abc$9276$new_n2536 ;
  wire \$abc$9276$new_n2537 ;
  wire \$abc$9276$new_n2538 ;
  wire \$abc$9276$new_n2539 ;
  wire \$abc$9276$new_n2540 ;
  wire \$abc$9276$new_n2541 ;
  wire \$abc$9276$new_n2542 ;
  wire \$abc$9276$new_n2543 ;
  wire \$abc$9276$new_n2544 ;
  wire \$abc$9276$new_n2545 ;
  wire \$abc$9276$new_n2546 ;
  wire \$abc$9276$new_n2547 ;
  wire \$abc$9276$new_n2548 ;
  wire \$abc$9276$new_n2549 ;
  wire \$abc$9276$new_n2550 ;
  wire \$abc$9276$new_n2551 ;
  wire \$abc$9276$new_n2552 ;
  wire \$abc$9276$new_n2553 ;
  wire \$abc$9276$new_n2554 ;
  wire \$abc$9276$new_n2555 ;
  wire \$abc$9276$new_n2556 ;
  wire \$abc$9276$new_n2557 ;
  wire \$abc$9276$new_n2558 ;
  wire \$abc$9276$new_n2559 ;
  wire \$abc$9276$new_n2560 ;
  wire \$abc$9276$new_n2561 ;
  wire \$abc$9276$new_n2562 ;
  wire \$abc$9276$new_n2563 ;
  wire \$abc$9276$new_n2564 ;
  wire \$abc$9276$new_n2565 ;
  wire \$abc$9276$new_n2566 ;
  wire \$abc$9276$new_n2567 ;
  wire \$abc$9276$new_n2568 ;
  wire \$abc$9276$new_n2569 ;
  wire \$abc$9276$new_n2570 ;
  wire \$abc$9276$new_n2571 ;
  wire \$abc$9276$new_n2572 ;
  wire \$abc$9276$new_n2573 ;
  wire \$abc$9276$new_n2575 ;
  wire \$abc$9276$new_n2576 ;
  wire \$abc$9276$new_n2578 ;
  wire \$abc$9276$new_n2579 ;
  wire \$abc$9276$new_n2580 ;
  wire \$abc$9276$new_n2581 ;
  wire \$abc$9276$new_n2582 ;
  wire \$abc$9276$new_n2584 ;
  wire \$abc$9276$new_n2585 ;
  wire \$abc$9276$new_n2586 ;
  wire \$abc$9276$new_n2588 ;
  wire \$abc$9276$new_n2589 ;
  wire \$abc$9276$new_n2590 ;
  wire \$abc$9276$new_n2592 ;
  wire \$abc$9276$new_n2593 ;
  wire \$abc$9276$new_n2594 ;
  wire \$abc$9276$new_n2596 ;
  wire \$abc$9276$new_n2597 ;
  wire \$abc$9276$new_n2598 ;
  wire \$abc$9276$new_n2599 ;
  wire \$abc$9276$new_n2600 ;
  wire \$abc$9276$new_n2602 ;
  wire \$abc$9276$new_n2603 ;
  wire \$abc$9276$new_n2604 ;
  wire \$abc$9276$new_n2605 ;
  wire \$abc$9276$new_n2606 ;
  wire \$abc$9276$new_n2608 ;
  wire \$abc$9276$new_n2609 ;
  wire \$abc$9276$new_n2610 ;
  wire \$abc$9276$new_n2611 ;
  wire \$abc$9276$new_n2612 ;
  wire \$abc$9276$new_n2614 ;
  wire \$abc$9276$new_n2615 ;
  wire \$abc$9276$new_n2617 ;
  wire \$abc$9276$new_n2618 ;
  wire \$abc$9276$new_n2619 ;
  wire \$abc$9276$new_n2620 ;
  wire \$abc$9276$new_n2621 ;
  wire \$abc$9276$new_n2622 ;
  wire \$abc$9276$new_n2623 ;
  wire \$abc$9276$new_n2624 ;
  wire \$abc$9276$new_n2625 ;
  wire \$abc$9276$new_n2626 ;
  wire \$abc$9276$new_n2627 ;
  wire \$abc$9276$new_n2628 ;
  wire \$abc$9276$new_n2629 ;
  wire \$abc$9276$new_n2630 ;
  wire \$abc$9276$new_n2631 ;
  wire \$abc$9276$new_n2633 ;
  wire \$abc$9276$new_n2634 ;
  wire \$abc$9276$new_n2635 ;
  wire \$abc$9276$new_n2636 ;
  wire \$abc$9276$new_n2637 ;
  wire \$abc$9276$new_n2638 ;
  wire \$abc$9276$new_n2640 ;
  wire \$abc$9276$new_n2641 ;
  wire \$abc$9276$new_n2642 ;
  wire \$abc$9276$new_n2643 ;
  wire \$abc$9276$new_n2645 ;
  wire \$abc$9276$new_n2646 ;
  wire \$abc$9276$new_n2647 ;
  wire \$abc$9276$new_n2648 ;
  wire \$abc$9276$new_n2649 ;
  wire \$abc$9276$new_n2650 ;
  wire \$abc$9276$new_n2651 ;
  wire \$abc$9276$new_n2652 ;
  wire \$abc$9276$new_n2654 ;
  wire \$abc$9276$new_n2655 ;
  wire \$abc$9276$new_n2656 ;
  wire \$abc$9276$new_n2657 ;
  wire \$abc$9276$new_n2658 ;
  wire \$abc$9276$new_n2659 ;
  wire \$abc$9276$new_n2660 ;
  wire \$abc$9276$new_n2661 ;
  wire \$abc$9276$new_n2662 ;
  wire \$abc$9276$new_n2663 ;
  wire \$abc$9276$new_n2664 ;
  wire \$abc$9276$new_n2665 ;
  wire \$abc$9276$new_n2666 ;
  wire \$abc$9276$new_n2667 ;
  wire \$abc$9276$new_n2668 ;
  wire \$abc$9276$new_n2669 ;
  wire \$abc$9276$new_n2671 ;
  wire \$abc$9276$new_n2672 ;
  wire \$abc$9276$new_n2673 ;
  wire \$abc$9276$new_n2674 ;
  wire \$abc$9276$new_n2675 ;
  wire \$abc$9276$new_n2676 ;
  wire \$abc$9276$new_n2678 ;
  wire \$abc$9276$new_n2679 ;
  wire \$abc$9276$new_n2680 ;
  wire \$abc$9276$new_n2681 ;
  wire \$abc$9276$new_n2682 ;
  wire \$abc$9276$new_n2683 ;
  wire \$abc$9276$new_n2684 ;
  wire \$abc$9276$new_n2685 ;
  wire \$abc$9276$new_n2686 ;
  wire \$abc$9276$new_n2687 ;
  wire \$abc$9276$new_n2688 ;
  wire \$abc$9276$new_n2689 ;
  wire \$abc$9276$new_n2690 ;
  wire \$abc$9276$new_n2691 ;
  wire \$abc$9276$new_n2693 ;
  wire \$abc$9276$new_n2694 ;
  wire \$abc$9276$new_n2695 ;
  wire \$abc$9276$new_n2696 ;
  wire \$abc$9276$new_n2697 ;
  wire \$abc$9276$new_n2698 ;
  wire \$abc$9276$new_n2699 ;
  wire \$abc$9276$new_n2700 ;
  wire \$abc$9276$new_n2701 ;
  wire \$abc$9276$new_n2702 ;
  wire \$abc$9276$new_n2703 ;
  wire \$abc$9276$new_n2705 ;
  wire \$abc$9276$new_n2706 ;
  wire \$abc$9276$new_n2707 ;
  wire \$abc$9276$new_n2708 ;
  wire \$abc$9276$new_n2709 ;
  wire \$abc$9276$new_n2710 ;
  wire \$abc$9276$new_n2711 ;
  wire \$abc$9276$new_n2712 ;
  wire \$abc$9276$new_n2713 ;
  wire \$abc$9276$new_n2714 ;
  wire \$abc$9276$new_n2715 ;
  wire \$abc$9276$new_n2717 ;
  wire \$abc$9276$new_n2718 ;
  wire \$abc$9276$new_n2719 ;
  wire \$abc$9276$new_n2720 ;
  wire \$abc$9276$new_n2721 ;
  wire \$abc$9276$new_n2722 ;
  wire \$abc$9276$new_n2723 ;
  wire \$abc$9276$new_n2724 ;
  wire \$abc$9276$new_n2725 ;
  wire \$abc$9276$new_n2727 ;
  wire \$abc$9276$new_n2728 ;
  wire \$abc$9276$new_n2729 ;
  wire \$abc$9276$new_n2730 ;
  wire \$abc$9276$new_n2731 ;
  wire \$abc$9276$new_n2732 ;
  wire \$abc$9276$new_n2733 ;
  wire \$abc$9276$new_n2734 ;
  wire \$abc$9276$new_n2735 ;
  wire \$abc$9276$new_n2736 ;
  wire \$abc$9276$new_n2737 ;
  wire \$abc$9276$new_n2738 ;
  wire \$abc$9276$new_n2740 ;
  wire \$abc$9276$new_n2741 ;
  wire \$abc$9276$new_n2742 ;
  wire \$abc$9276$new_n2743 ;
  wire \$abc$9276$new_n2744 ;
  wire \$abc$9276$new_n2745 ;
  wire \$abc$9276$new_n2746 ;
  wire \$abc$9276$new_n2747 ;
  wire \$abc$9276$new_n2748 ;
  wire \$abc$9276$new_n2749 ;
  wire \$abc$9276$new_n2751 ;
  wire \$abc$9276$new_n2752 ;
  wire \$abc$9276$new_n2753 ;
  wire \$abc$9276$new_n2754 ;
  wire \$abc$9276$new_n2755 ;
  wire \$abc$9276$new_n2756 ;
  wire \$abc$9276$new_n2757 ;
  wire \$abc$9276$new_n2758 ;
  wire \$abc$9276$new_n2759 ;
  wire \$abc$9276$new_n2760 ;
  wire \$abc$9276$new_n2761 ;
  wire \$abc$9276$new_n2763 ;
  wire \$abc$9276$new_n2764 ;
  wire \$abc$9276$new_n2765 ;
  wire \$abc$9276$new_n2766 ;
  wire \$abc$9276$new_n2767 ;
  wire \$abc$9276$new_n2768 ;
  wire \$abc$9276$new_n2769 ;
  wire \$abc$9276$new_n2770 ;
  wire \$abc$9276$new_n2771 ;
  wire \$abc$9276$new_n2772 ;
  wire \$abc$9276$new_n2773 ;
  wire \$abc$9276$new_n2775 ;
  wire \$abc$9276$new_n346 ;
  wire \$abc$9276$new_n347 ;
  wire \$abc$9276$new_n348 ;
  wire \$abc$9276$new_n349 ;
  wire \$abc$9276$new_n350 ;
  wire \$abc$9276$new_n351 ;
  wire \$abc$9276$new_n352 ;
  wire \$abc$9276$new_n353 ;
  wire \$abc$9276$new_n354 ;
  wire \$abc$9276$new_n355 ;
  wire \$abc$9276$new_n356 ;
  wire \$abc$9276$new_n357 ;
  wire \$abc$9276$new_n358 ;
  wire \$abc$9276$new_n359 ;
  wire \$abc$9276$new_n360 ;
  wire \$abc$9276$new_n361 ;
  wire \$abc$9276$new_n362 ;
  wire \$abc$9276$new_n363 ;
  wire \$abc$9276$new_n364 ;
  wire \$abc$9276$new_n365 ;
  wire \$abc$9276$new_n366 ;
  wire \$abc$9276$new_n367 ;
  wire \$abc$9276$new_n368 ;
  wire \$abc$9276$new_n369 ;
  wire \$abc$9276$new_n370 ;
  wire \$abc$9276$new_n371 ;
  wire \$abc$9276$new_n372 ;
  wire \$abc$9276$new_n373 ;
  wire \$abc$9276$new_n374 ;
  wire \$abc$9276$new_n375 ;
  wire \$abc$9276$new_n376 ;
  wire \$abc$9276$new_n377 ;
  wire \$abc$9276$new_n378 ;
  wire \$abc$9276$new_n379 ;
  wire \$abc$9276$new_n380 ;
  wire \$abc$9276$new_n381 ;
  wire \$abc$9276$new_n382 ;
  wire \$abc$9276$new_n383 ;
  wire \$abc$9276$new_n384 ;
  wire \$abc$9276$new_n385 ;
  wire \$abc$9276$new_n386 ;
  wire \$abc$9276$new_n387 ;
  wire \$abc$9276$new_n388 ;
  wire \$abc$9276$new_n389 ;
  wire \$abc$9276$new_n390 ;
  wire \$abc$9276$new_n391 ;
  wire \$abc$9276$new_n392 ;
  wire \$abc$9276$new_n393 ;
  wire \$abc$9276$new_n394 ;
  wire \$abc$9276$new_n395 ;
  wire \$abc$9276$new_n396 ;
  wire \$abc$9276$new_n397 ;
  wire \$abc$9276$new_n398 ;
  wire \$abc$9276$new_n399 ;
  wire \$abc$9276$new_n400 ;
  wire \$abc$9276$new_n401 ;
  wire \$abc$9276$new_n402 ;
  wire \$abc$9276$new_n403 ;
  wire \$abc$9276$new_n404 ;
  wire \$abc$9276$new_n405 ;
  wire \$abc$9276$new_n406 ;
  wire \$abc$9276$new_n407 ;
  wire \$abc$9276$new_n408 ;
  wire \$abc$9276$new_n409 ;
  wire \$abc$9276$new_n410 ;
  wire \$abc$9276$new_n411 ;
  wire \$abc$9276$new_n412 ;
  wire \$abc$9276$new_n413 ;
  wire \$abc$9276$new_n414 ;
  wire \$abc$9276$new_n415 ;
  wire \$abc$9276$new_n416 ;
  wire \$abc$9276$new_n417 ;
  wire \$abc$9276$new_n418 ;
  wire \$abc$9276$new_n419 ;
  wire \$abc$9276$new_n420 ;
  wire \$abc$9276$new_n421 ;
  wire \$abc$9276$new_n422 ;
  wire \$abc$9276$new_n423 ;
  wire \$abc$9276$new_n424 ;
  wire \$abc$9276$new_n425 ;
  wire \$abc$9276$new_n426 ;
  wire \$abc$9276$new_n427 ;
  wire \$abc$9276$new_n428 ;
  wire \$abc$9276$new_n429 ;
  wire \$abc$9276$new_n430 ;
  wire \$abc$9276$new_n431 ;
  wire \$abc$9276$new_n432 ;
  wire \$abc$9276$new_n433 ;
  wire \$abc$9276$new_n434 ;
  wire \$abc$9276$new_n435 ;
  wire \$abc$9276$new_n436 ;
  wire \$abc$9276$new_n437 ;
  wire \$abc$9276$new_n438 ;
  wire \$abc$9276$new_n439 ;
  wire \$abc$9276$new_n440 ;
  wire \$abc$9276$new_n441 ;
  wire \$abc$9276$new_n442 ;
  wire \$abc$9276$new_n443 ;
  wire \$abc$9276$new_n444 ;
  wire \$abc$9276$new_n445 ;
  wire \$abc$9276$new_n446 ;
  wire \$abc$9276$new_n447 ;
  wire \$abc$9276$new_n448 ;
  wire \$abc$9276$new_n449 ;
  wire \$abc$9276$new_n450 ;
  wire \$abc$9276$new_n451 ;
  wire \$abc$9276$new_n452 ;
  wire \$abc$9276$new_n453 ;
  wire \$abc$9276$new_n454 ;
  wire \$abc$9276$new_n455 ;
  wire \$abc$9276$new_n456 ;
  wire \$abc$9276$new_n457 ;
  wire \$abc$9276$new_n458 ;
  wire \$abc$9276$new_n459 ;
  wire \$abc$9276$new_n460 ;
  wire \$abc$9276$new_n461 ;
  wire \$abc$9276$new_n462 ;
  wire \$abc$9276$new_n463 ;
  wire \$abc$9276$new_n464 ;
  wire \$abc$9276$new_n465 ;
  wire \$abc$9276$new_n466 ;
  wire \$abc$9276$new_n467 ;
  wire \$abc$9276$new_n468 ;
  wire \$abc$9276$new_n469 ;
  wire \$abc$9276$new_n470 ;
  wire \$abc$9276$new_n471 ;
  wire \$abc$9276$new_n472 ;
  wire \$abc$9276$new_n473 ;
  wire \$abc$9276$new_n474 ;
  wire \$abc$9276$new_n475 ;
  wire \$abc$9276$new_n476 ;
  wire \$abc$9276$new_n477 ;
  wire \$abc$9276$new_n478 ;
  wire \$abc$9276$new_n479 ;
  wire \$abc$9276$new_n480 ;
  wire \$abc$9276$new_n481 ;
  wire \$abc$9276$new_n482 ;
  wire \$abc$9276$new_n483 ;
  wire \$abc$9276$new_n484 ;
  wire \$abc$9276$new_n485 ;
  wire \$abc$9276$new_n486 ;
  wire \$abc$9276$new_n487 ;
  wire \$abc$9276$new_n489 ;
  wire \$abc$9276$new_n490 ;
  wire \$abc$9276$new_n491 ;
  wire \$abc$9276$new_n492 ;
  wire \$abc$9276$new_n493 ;
  wire \$abc$9276$new_n494 ;
  wire \$abc$9276$new_n496 ;
  wire \$abc$9276$new_n497 ;
  wire \$abc$9276$new_n498 ;
  wire \$abc$9276$new_n499 ;
  wire \$abc$9276$new_n500 ;
  wire \$abc$9276$new_n501 ;
  wire \$abc$9276$new_n502 ;
  wire \$abc$9276$new_n503 ;
  wire \$abc$9276$new_n504 ;
  wire \$abc$9276$new_n505 ;
  wire \$abc$9276$new_n507 ;
  wire \$abc$9276$new_n508 ;
  wire \$abc$9276$new_n509 ;
  wire \$abc$9276$new_n510 ;
  wire \$abc$9276$new_n511 ;
  wire \$abc$9276$new_n512 ;
  wire \$abc$9276$new_n514 ;
  wire \$abc$9276$new_n515 ;
  wire \$abc$9276$new_n516 ;
  wire \$abc$9276$new_n517 ;
  wire \$abc$9276$new_n518 ;
  wire \$abc$9276$new_n519 ;
  wire \$abc$9276$new_n520 ;
  wire \$abc$9276$new_n521 ;
  wire \$abc$9276$new_n522 ;
  wire \$abc$9276$new_n523 ;
  wire \$abc$9276$new_n524 ;
  wire \$abc$9276$new_n525 ;
  wire \$abc$9276$new_n527 ;
  wire \$abc$9276$new_n528 ;
  wire \$abc$9276$new_n529 ;
  wire \$abc$9276$new_n530 ;
  wire \$abc$9276$new_n531 ;
  wire \$abc$9276$new_n532 ;
  wire \$abc$9276$new_n534 ;
  wire \$abc$9276$new_n535 ;
  wire \$abc$9276$new_n536 ;
  wire \$abc$9276$new_n537 ;
  wire \$abc$9276$new_n538 ;
  wire \$abc$9276$new_n539 ;
  wire \$abc$9276$new_n540 ;
  wire \$abc$9276$new_n541 ;
  wire \$abc$9276$new_n542 ;
  wire \$abc$9276$new_n543 ;
  wire \$abc$9276$new_n544 ;
  wire \$abc$9276$new_n545 ;
  wire \$abc$9276$new_n547 ;
  wire \$abc$9276$new_n548 ;
  wire \$abc$9276$new_n549 ;
  wire \$abc$9276$new_n550 ;
  wire \$abc$9276$new_n551 ;
  wire \$abc$9276$new_n552 ;
  wire \$abc$9276$new_n554 ;
  wire \$abc$9276$new_n555 ;
  wire \$abc$9276$new_n556 ;
  wire \$abc$9276$new_n557 ;
  wire \$abc$9276$new_n558 ;
  wire \$abc$9276$new_n559 ;
  wire \$abc$9276$new_n560 ;
  wire \$abc$9276$new_n561 ;
  wire \$abc$9276$new_n562 ;
  wire \$abc$9276$new_n563 ;
  wire \$abc$9276$new_n564 ;
  wire \$abc$9276$new_n565 ;
  wire \$abc$9276$new_n566 ;
  wire \$abc$9276$new_n567 ;
  wire \$abc$9276$new_n568 ;
  wire \$abc$9276$new_n570 ;
  wire \$abc$9276$new_n571 ;
  wire \$abc$9276$new_n572 ;
  wire \$abc$9276$new_n573 ;
  wire \$abc$9276$new_n574 ;
  wire \$abc$9276$new_n575 ;
  wire \$abc$9276$new_n577 ;
  wire \$abc$9276$new_n578 ;
  wire \$abc$9276$new_n579 ;
  wire \$abc$9276$new_n580 ;
  wire \$abc$9276$new_n581 ;
  wire \$abc$9276$new_n582 ;
  wire \$abc$9276$new_n583 ;
  wire \$abc$9276$new_n584 ;
  wire \$abc$9276$new_n585 ;
  wire \$abc$9276$new_n586 ;
  wire \$abc$9276$new_n588 ;
  wire \$abc$9276$new_n589 ;
  wire \$abc$9276$new_n590 ;
  wire \$abc$9276$new_n591 ;
  wire \$abc$9276$new_n592 ;
  wire \$abc$9276$new_n593 ;
  wire \$abc$9276$new_n595 ;
  wire \$abc$9276$new_n596 ;
  wire \$abc$9276$new_n597 ;
  wire \$abc$9276$new_n598 ;
  wire \$abc$9276$new_n599 ;
  wire \$abc$9276$new_n600 ;
  wire \$abc$9276$new_n601 ;
  wire \$abc$9276$new_n602 ;
  wire \$abc$9276$new_n603 ;
  wire \$abc$9276$new_n604 ;
  wire \$abc$9276$new_n605 ;
  wire \$abc$9276$new_n606 ;
  wire \$abc$9276$new_n608 ;
  wire \$abc$9276$new_n609 ;
  wire \$abc$9276$new_n610 ;
  wire \$abc$9276$new_n611 ;
  wire \$abc$9276$new_n612 ;
  wire \$abc$9276$new_n613 ;
  wire \$abc$9276$new_n615 ;
  wire \$abc$9276$new_n616 ;
  wire \$abc$9276$new_n617 ;
  wire \$abc$9276$new_n618 ;
  wire \$abc$9276$new_n619 ;
  wire \$abc$9276$new_n620 ;
  wire \$abc$9276$new_n621 ;
  wire \$abc$9276$new_n622 ;
  wire \$abc$9276$new_n623 ;
  wire \$abc$9276$new_n624 ;
  wire \$abc$9276$new_n626 ;
  wire \$abc$9276$new_n627 ;
  wire \$abc$9276$new_n628 ;
  wire \$abc$9276$new_n629 ;
  wire \$abc$9276$new_n630 ;
  wire \$abc$9276$new_n631 ;
  wire \$abc$9276$new_n633 ;
  wire \$abc$9276$new_n634 ;
  wire \$abc$9276$new_n635 ;
  wire \$abc$9276$new_n637 ;
  wire \$abc$9276$new_n638 ;
  wire \$abc$9276$new_n640 ;
  wire \$abc$9276$new_n641 ;
  wire \$abc$9276$new_n643 ;
  wire \$abc$9276$new_n644 ;
  wire \$abc$9276$new_n646 ;
  wire \$abc$9276$new_n647 ;
  wire \$abc$9276$new_n649 ;
  wire \$abc$9276$new_n650 ;
  wire \$abc$9276$new_n652 ;
  wire \$abc$9276$new_n653 ;
  wire \$abc$9276$new_n655 ;
  wire \$abc$9276$new_n656 ;
  wire \$abc$9276$new_n658 ;
  wire \$abc$9276$new_n659 ;
  wire \$abc$9276$new_n660 ;
  wire \$abc$9276$new_n661 ;
  wire \$abc$9276$new_n663 ;
  wire \$abc$9276$new_n664 ;
  wire \$abc$9276$new_n666 ;
  wire \$abc$9276$new_n667 ;
  wire \$abc$9276$new_n669 ;
  wire \$abc$9276$new_n670 ;
  wire \$abc$9276$new_n672 ;
  wire \$abc$9276$new_n673 ;
  wire \$abc$9276$new_n675 ;
  wire \$abc$9276$new_n676 ;
  wire \$abc$9276$new_n678 ;
  wire \$abc$9276$new_n679 ;
  wire \$abc$9276$new_n681 ;
  wire \$abc$9276$new_n682 ;
  wire \$abc$9276$new_n684 ;
  wire \$abc$9276$new_n685 ;
  wire \$abc$9276$new_n686 ;
  wire \$abc$9276$new_n687 ;
  wire \$abc$9276$new_n689 ;
  wire \$abc$9276$new_n690 ;
  wire \$abc$9276$new_n692 ;
  wire \$abc$9276$new_n693 ;
  wire \$abc$9276$new_n695 ;
  wire \$abc$9276$new_n696 ;
  wire \$abc$9276$new_n698 ;
  wire \$abc$9276$new_n699 ;
  wire \$abc$9276$new_n701 ;
  wire \$abc$9276$new_n702 ;
  wire \$abc$9276$new_n704 ;
  wire \$abc$9276$new_n705 ;
  wire \$abc$9276$new_n707 ;
  wire \$abc$9276$new_n708 ;
  wire \$abc$9276$new_n710 ;
  wire \$abc$9276$new_n711 ;
  wire \$abc$9276$new_n712 ;
  wire \$abc$9276$new_n713 ;
  wire \$abc$9276$new_n714 ;
  wire \$abc$9276$new_n715 ;
  wire \$abc$9276$new_n716 ;
  wire \$abc$9276$new_n717 ;
  wire \$abc$9276$new_n718 ;
  wire \$abc$9276$new_n719 ;
  wire \$abc$9276$new_n720 ;
  wire \$abc$9276$new_n721 ;
  wire \$abc$9276$new_n722 ;
  wire \$abc$9276$new_n723 ;
  wire \$abc$9276$new_n724 ;
  wire \$abc$9276$new_n725 ;
  wire \$abc$9276$new_n726 ;
  wire \$abc$9276$new_n727 ;
  wire \$abc$9276$new_n728 ;
  wire \$abc$9276$new_n729 ;
  wire \$abc$9276$new_n730 ;
  wire \$abc$9276$new_n731 ;
  wire \$abc$9276$new_n732 ;
  wire \$abc$9276$new_n733 ;
  wire \$abc$9276$new_n734 ;
  wire \$abc$9276$new_n735 ;
  wire \$abc$9276$new_n736 ;
  wire \$abc$9276$new_n737 ;
  wire \$abc$9276$new_n738 ;
  wire \$abc$9276$new_n739 ;
  wire \$abc$9276$new_n740 ;
  wire \$abc$9276$new_n741 ;
  wire \$abc$9276$new_n742 ;
  wire \$abc$9276$new_n743 ;
  wire \$abc$9276$new_n744 ;
  wire \$abc$9276$new_n745 ;
  wire \$abc$9276$new_n746 ;
  wire \$abc$9276$new_n747 ;
  wire \$abc$9276$new_n748 ;
  wire \$abc$9276$new_n749 ;
  wire \$abc$9276$new_n750 ;
  wire \$abc$9276$new_n752 ;
  wire \$abc$9276$new_n753 ;
  wire \$abc$9276$new_n754 ;
  wire \$abc$9276$new_n755 ;
  wire \$abc$9276$new_n756 ;
  wire \$abc$9276$new_n757 ;
  wire \$abc$9276$new_n758 ;
  wire \$abc$9276$new_n759 ;
  wire \$abc$9276$new_n760 ;
  wire \$abc$9276$new_n761 ;
  wire \$abc$9276$new_n762 ;
  wire \$abc$9276$new_n763 ;
  wire \$abc$9276$new_n764 ;
  wire \$abc$9276$new_n765 ;
  wire \$abc$9276$new_n766 ;
  wire \$abc$9276$new_n767 ;
  wire \$abc$9276$new_n768 ;
  wire \$abc$9276$new_n769 ;
  wire \$abc$9276$new_n770 ;
  wire \$abc$9276$new_n771 ;
  wire \$abc$9276$new_n772 ;
  wire \$abc$9276$new_n773 ;
  wire \$abc$9276$new_n774 ;
  wire \$abc$9276$new_n775 ;
  wire \$abc$9276$new_n776 ;
  wire \$abc$9276$new_n777 ;
  wire \$abc$9276$new_n778 ;
  wire \$abc$9276$new_n779 ;
  wire \$abc$9276$new_n780 ;
  wire \$abc$9276$new_n781 ;
  wire \$abc$9276$new_n782 ;
  wire \$abc$9276$new_n783 ;
  wire \$abc$9276$new_n784 ;
  wire \$abc$9276$new_n785 ;
  wire \$abc$9276$new_n786 ;
  wire \$abc$9276$new_n787 ;
  wire \$abc$9276$new_n788 ;
  wire \$abc$9276$new_n789 ;
  wire \$abc$9276$new_n790 ;
  wire \$abc$9276$new_n791 ;
  wire \$abc$9276$new_n792 ;
  wire \$abc$9276$new_n793 ;
  wire \$abc$9276$new_n794 ;
  wire \$abc$9276$new_n795 ;
  wire \$abc$9276$new_n796 ;
  wire \$abc$9276$new_n797 ;
  wire \$abc$9276$new_n798 ;
  wire \$abc$9276$new_n799 ;
  wire \$abc$9276$new_n800 ;
  wire \$abc$9276$new_n801 ;
  wire \$abc$9276$new_n802 ;
  wire \$abc$9276$new_n803 ;
  wire \$abc$9276$new_n804 ;
  wire \$abc$9276$new_n805 ;
  wire \$abc$9276$new_n806 ;
  wire \$abc$9276$new_n807 ;
  wire \$abc$9276$new_n808 ;
  wire \$abc$9276$new_n809 ;
  wire \$abc$9276$new_n810 ;
  wire \$abc$9276$new_n811 ;
  wire \$abc$9276$new_n812 ;
  wire \$abc$9276$new_n813 ;
  wire \$abc$9276$new_n814 ;
  wire \$abc$9276$new_n815 ;
  wire \$abc$9276$new_n816 ;
  wire \$abc$9276$new_n817 ;
  wire \$abc$9276$new_n818 ;
  wire \$abc$9276$new_n820 ;
  wire \$abc$9276$new_n821 ;
  wire \$abc$9276$new_n822 ;
  wire \$abc$9276$new_n823 ;
  wire \$abc$9276$new_n825 ;
  wire \$abc$9276$new_n826 ;
  wire \$abc$9276$new_n827 ;
  wire \$abc$9276$new_n828 ;
  wire \$abc$9276$new_n829 ;
  wire \$abc$9276$new_n830 ;
  wire \$abc$9276$new_n831 ;
  wire \$abc$9276$new_n833 ;
  wire \$abc$9276$new_n834 ;
  wire \$abc$9276$new_n835 ;
  wire \$abc$9276$new_n836 ;
  wire \$abc$9276$new_n838 ;
  wire \$abc$9276$new_n839 ;
  wire \$abc$9276$new_n840 ;
  wire \$abc$9276$new_n842 ;
  wire \$abc$9276$new_n843 ;
  wire \$abc$9276$new_n845 ;
  wire \$abc$9276$new_n846 ;
  wire \$abc$9276$new_n847 ;
  wire \$abc$9276$new_n849 ;
  wire \$abc$9276$new_n850 ;
  wire \$abc$9276$new_n852 ;
  wire \$abc$9276$new_n853 ;
  wire \$abc$9276$new_n854 ;
  wire \$abc$9276$new_n855 ;
  wire \$abc$9276$new_n857 ;
  wire \$abc$9276$new_n858 ;
  wire \$abc$9276$new_n859 ;
  wire \$abc$9276$new_n860 ;
  wire \$abc$9276$new_n861 ;
  wire \$abc$9276$new_n863 ;
  wire \$abc$9276$new_n864 ;
  wire \$abc$9276$new_n865 ;
  wire \$abc$9276$new_n866 ;
  wire \$abc$9276$new_n867 ;
  wire \$abc$9276$new_n868 ;
  wire \$abc$9276$new_n869 ;
  wire \$abc$9276$new_n870 ;
  wire \$abc$9276$new_n871 ;
  wire \$abc$9276$new_n872 ;
  wire \$abc$9276$new_n874 ;
  wire \$abc$9276$new_n875 ;
  wire \$abc$9276$new_n876 ;
  wire \$abc$9276$new_n878 ;
  wire \$abc$9276$new_n879 ;
  wire \$abc$9276$new_n880 ;
  wire \$abc$9276$new_n881 ;
  wire \$abc$9276$new_n882 ;
  wire \$abc$9276$new_n883 ;
  wire \$abc$9276$new_n884 ;
  wire \$abc$9276$new_n885 ;
  wire \$abc$9276$new_n886 ;
  wire \$abc$9276$new_n887 ;
  wire \$abc$9276$new_n888 ;
  wire \$abc$9276$new_n889 ;
  wire \$abc$9276$new_n890 ;
  wire \$abc$9276$new_n891 ;
  wire \$abc$9276$new_n892 ;
  wire \$abc$9276$new_n893 ;
  wire \$abc$9276$new_n894 ;
  wire \$abc$9276$new_n895 ;
  wire \$abc$9276$new_n896 ;
  wire \$abc$9276$new_n898 ;
  wire \$abc$9276$new_n900 ;
  wire \$abc$9276$new_n901 ;
  wire \$abc$9276$new_n902 ;
  wire \$abc$9276$new_n903 ;
  wire \$abc$9276$new_n904 ;
  wire \$abc$9276$new_n905 ;
  wire \$abc$9276$new_n907 ;
  wire \$abc$9276$new_n908 ;
  wire \$abc$9276$new_n909 ;
  wire \$abc$9276$new_n911 ;
  wire \$abc$9276$new_n912 ;
  wire \$abc$9276$new_n913 ;
  wire \$abc$9276$new_n914 ;
  wire \$abc$9276$new_n915 ;
  wire \$abc$9276$new_n916 ;
  wire \$abc$9276$new_n918 ;
  wire \$abc$9276$new_n919 ;
  wire \$abc$9276$new_n920 ;
  wire \$abc$9276$new_n922 ;
  wire \$abc$9276$new_n923 ;
  wire \$abc$9276$new_n924 ;
  wire \$abc$9276$new_n926 ;
  wire \$abc$9276$new_n927 ;
  wire \$abc$9276$new_n928 ;
  wire \$abc$9276$new_n929 ;
  wire \$abc$9276$new_n930 ;
  wire \$abc$9276$new_n932 ;
  wire \$abc$9276$new_n933 ;
  wire \$abc$9276$new_n934 ;
  wire \$abc$9276$new_n935 ;
  wire \$abc$9276$new_n936 ;
  wire \$abc$9276$new_n937 ;
  wire \$abc$9276$new_n938 ;
  wire \$abc$9276$new_n939 ;
  wire \$abc$9276$new_n940 ;
  wire \$abc$9276$new_n941 ;
  wire \$abc$9276$new_n942 ;
  wire \$abc$9276$new_n943 ;
  wire \$abc$9276$new_n944 ;
  wire \$abc$9276$new_n946 ;
  wire \$abc$9276$new_n947 ;
  wire \$abc$9276$new_n948 ;
  wire \$abc$9276$new_n949 ;
  wire \$abc$9276$new_n950 ;
  wire \$abc$9276$new_n951 ;
  wire \$abc$9276$new_n952 ;
  wire \$abc$9276$new_n953 ;
  wire \$abc$9276$new_n954 ;
  wire \$abc$9276$new_n955 ;
  wire \$abc$9276$new_n956 ;
  wire \$abc$9276$new_n957 ;
  wire \$abc$9276$new_n958 ;
  wire \$abc$9276$new_n959 ;
  wire \$abc$9276$new_n960 ;
  wire \$abc$9276$new_n961 ;
  wire \$abc$9276$new_n962 ;
  wire \$abc$9276$new_n963 ;
  wire \$abc$9276$new_n964 ;
  wire \$abc$9276$new_n965 ;
  wire \$abc$9276$new_n966 ;
  wire \$abc$9276$new_n967 ;
  wire \$abc$9276$new_n968 ;
  wire \$abc$9276$new_n969 ;
  wire \$abc$9276$new_n970 ;
  wire \$abc$9276$new_n971 ;
  wire \$abc$9276$new_n972 ;
  wire \$abc$9276$new_n973 ;
  wire \$abc$9276$new_n975 ;
  wire \$abc$9276$new_n976 ;
  wire \$abc$9276$new_n977 ;
  wire \$abc$9276$new_n978 ;
  wire \$abc$9276$new_n979 ;
  wire \$abc$9276$new_n980 ;
  wire \$abc$9276$new_n981 ;
  wire \$abc$9276$new_n982 ;
  wire \$abc$9276$new_n983 ;
  wire \$abc$9276$new_n984 ;
  wire \$abc$9276$new_n985 ;
  wire \$abc$9276$new_n986 ;
  wire \$abc$9276$new_n987 ;
  wire \$abc$9276$new_n988 ;
  wire \$abc$9276$new_n989 ;
  wire \$abc$9276$new_n990 ;
  wire \$abc$9276$new_n991 ;
  wire \$abc$9276$new_n992 ;
  wire \$abc$9276$new_n993 ;
  wire \$abc$9276$new_n994 ;
  wire \$abc$9276$new_n995 ;
  wire \$abc$9276$new_n996 ;
  wire \$abc$9276$new_n997 ;
  wire \$abc$9276$new_n998 ;
  wire \$abc$9276$new_n999 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9112 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9113 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9114 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9115 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9116 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9117 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9118 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9119 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9122 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9123 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9124 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9125 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9126 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9127 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9128 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9129 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9130 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9131 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9144 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9145 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9146 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9147 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9148 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9149 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9150 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9151 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9152 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9153 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9154 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9155 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9156 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9157 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9158 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9159 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9162 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9163 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9164 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9165 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9166 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9167 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9168 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9169 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9178 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9179 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9186 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9187 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9188 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9189 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9190 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9191 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9192 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9193 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9194 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9195 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9196 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9197 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9198 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9199 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9200 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9201 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9202 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9203 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9204 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9205 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9208 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9209 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9212 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9213 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9214 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9215 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9216 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9217 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9218 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9219 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9220 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9221 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9222 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9223 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9224 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9225 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9232 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9233 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9234 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9235 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9236 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9237 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9238 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9239 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9240 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9241 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9242 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9243 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9244 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9245 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9246 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9247 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9248 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9249 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9250 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9251 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9252 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9253 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9254 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9255 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9256 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9257 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9258 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9259 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9260 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9261 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9262 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9263 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9268 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9269 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9270 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9271 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9272 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9273 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9274 ;
  wire \$auto$dfflibmap.cc:532:dfflibmap$9275 ;
  wire \$auto$hilomap.cc:39:hilomap_worker$12030 ;
  wire \$flatten \CPU.\$procmux$291.B ;
  wire \$flatten \CPU.\$procmux$415.B ;
  wire \$flatten \CPU.\$procmux$715.B ;
  wire CPU.ABH;
  wire CPU.ABL;
  wire CPU.ADD;
  wire CPU.ALU.AI7;
  wire CPU.ALU.BI7;
  wire CPU.ALU.CO;
  wire CPU.ALU.HC;
  wire CPU.ALU.N;
  wire CPU.AXYS[0];
  wire CPU.AXYS[1];
  wire CPU.AXYS[2];
  wire CPU.AXYS[3];
  wire CPU.C;
  wire CPU.D;
  wire CPU.DIHOLD;
  wire CPU.DIMUX;
  wire CPU.I;
  wire CPU.IRHOLD;
  wire CPU.IRHOLD_valid;
  wire CPU.N;
  wire CPU.NMI_1;
  wire CPU.NMI_edge;
  wire CPU.PC;
  wire CPU.V;
  wire CPU.Z;
  wire CPU.adc_bcd;
  wire CPU.adc_sbc;
  wire CPU.adj_bcd;
  wire CPU.backwards;
  wire CPU.bit_ins;
  wire CPU.clc;
  wire CPU.cld;
  wire CPU.cli;
  wire CPU.clv;
  wire CPU.compare;
  wire CPU.cond_code;
  wire CPU.dst_reg;
  wire CPU.inc;
  wire CPU.index_y;
  wire CPU.load_only;
  wire CPU.load_reg;
  wire CPU.op;
  wire CPU.php;
  wire CPU.plp;
  wire CPU.res;
  wire CPU.rotate;
  wire CPU.sec;
  wire CPU.sed;
  wire CPU.sei;
  wire CPU.shift;
  wire CPU.shift_right;
  wire CPU.src_reg;
  wire CPU.state;
  wire CPU.store;
  wire CPU.write_back;
  wire clk_cts_n0;
  wire clk_cts_n1;
  wire clk_cts_n2;
  wire clk_cts_n3;
  wire clk_cts_n4;
  wire clk_cts_n5;
  wire clk_cts_n6;
  wire clk_cts_n7;
  wire clk_cts_n8;
  wire clk_cts_n9;
  wire clk_cts_n10;
  wire clk_cts_n11;
  wire clk_cts_n12;
  wire clk_cts_n13;
  wire clk_cts_n14;
  wire clk_cts_n15;
  wire clk_cts_n16;
  wire clk_cts_n17;
  wire clk_cts_n18;
  wire clk_cts_n19;
  wire clk_cts_n20;
  wire clk_cts_n21;
  wire clk_cts_n22;
  wire clk_cts_n23;
  wire clk_cts_n24;
  wire clk_cts_n25;
  wire clk_cts_n26;
  wire clk_cts_n27;
  wire clk_cts_n28;
  wire clk_cts_n29;
  wire clk_cts_root;
  wire tie_low_T0Y0;
  wire tie_high_T0Y0;
  wire tie_low_T1Y0;
  wire tie_high_T1Y0;
  wire tie_low_T2Y0;
  wire tie_high_T2Y0;
  wire tie_low_T3Y0;
  wire tie_high_T3Y0;
  wire tie_low_T4Y0;
  wire tie_high_T4Y0;
  wire tie_low_T5Y0;
  wire tie_high_T5Y0;
  wire tie_low_T6Y0;
  wire tie_high_T6Y0;
  wire tie_low_T7Y0;
  wire tie_high_T7Y0;
  wire tie_low_T8Y0;
  wire tie_high_T8Y0;
  wire tie_low_T9Y0;
  wire tie_high_T9Y0;
  wire tie_low_T10Y0;
  wire tie_high_T10Y0;
  wire tie_low_T11Y0;
  wire tie_high_T11Y0;
  wire tie_low_T12Y0;
  wire tie_high_T12Y0;
  wire tie_low_T13Y0;
  wire tie_high_T13Y0;
  wire tie_low_T14Y0;
  wire tie_high_T14Y0;
  wire tie_low_T15Y0;
  wire tie_high_T15Y0;
  wire tie_low_T16Y0;
  wire tie_high_T16Y0;
  wire tie_low_T17Y0;
  wire tie_high_T17Y0;
  wire tie_low_T18Y0;
  wire tie_high_T18Y0;
  wire tie_low_T19Y0;
  wire tie_high_T19Y0;
  wire tie_low_T20Y0;
  wire tie_high_T20Y0;
  wire tie_low_T21Y0;
  wire tie_high_T21Y0;
  wire tie_low_T22Y0;
  wire tie_high_T22Y0;
  wire tie_low_T23Y0;
  wire tie_high_T23Y0;
  wire tie_low_T24Y0;
  wire tie_high_T24Y0;
  wire tie_low_T25Y0;
  wire tie_high_T25Y0;
  wire tie_low_T26Y0;
  wire tie_high_T26Y0;
  wire tie_low_T27Y0;
  wire tie_high_T27Y0;
  wire tie_low_T28Y0;
  wire tie_high_T28Y0;
  wire tie_low_T29Y0;
  wire tie_high_T29Y0;
  wire tie_low_T30Y0;
  wire tie_high_T30Y0;
  wire tie_low_T31Y0;
  wire tie_high_T31Y0;
  wire tie_low_T32Y0;
  wire tie_high_T32Y0;
  wire tie_low_T33Y0;
  wire tie_high_T33Y0;
  wire tie_low_T34Y0;
  wire tie_high_T34Y0;
  wire tie_low_T35Y0;
  wire tie_high_T35Y0;
  wire tie_low_T0Y1;
  wire tie_high_T0Y1;
  wire tie_low_T1Y1;
  wire tie_high_T1Y1;
  wire tie_low_T2Y1;
  wire tie_high_T2Y1;
  wire tie_low_T3Y1;
  wire tie_high_T3Y1;
  wire tie_low_T4Y1;
  wire tie_high_T4Y1;
  wire tie_low_T5Y1;
  wire tie_high_T5Y1;
  wire tie_low_T6Y1;
  wire tie_high_T6Y1;
  wire tie_low_T7Y1;
  wire tie_high_T7Y1;
  wire tie_low_T8Y1;
  wire tie_high_T8Y1;
  wire tie_low_T9Y1;
  wire tie_high_T9Y1;
  wire tie_low_T10Y1;
  wire tie_high_T10Y1;
  wire tie_low_T11Y1;
  wire tie_high_T11Y1;
  wire tie_low_T12Y1;
  wire tie_high_T12Y1;
  wire tie_low_T13Y1;
  wire tie_high_T13Y1;
  wire tie_low_T14Y1;
  wire tie_high_T14Y1;
  wire tie_low_T15Y1;
  wire tie_high_T15Y1;
  wire tie_low_T16Y1;
  wire tie_high_T16Y1;
  wire tie_low_T17Y1;
  wire tie_high_T17Y1;
  wire tie_low_T18Y1;
  wire tie_high_T18Y1;
  wire tie_low_T19Y1;
  wire tie_high_T19Y1;
  wire tie_low_T20Y1;
  wire tie_high_T20Y1;
  wire tie_low_T21Y1;
  wire tie_high_T21Y1;
  wire tie_low_T22Y1;
  wire tie_high_T22Y1;
  wire tie_low_T23Y1;
  wire tie_high_T23Y1;
  wire tie_low_T24Y1;
  wire tie_high_T24Y1;
  wire tie_low_T25Y1;
  wire tie_high_T25Y1;
  wire tie_low_T26Y1;
  wire tie_high_T26Y1;
  wire tie_low_T27Y1;
  wire tie_high_T27Y1;
  wire tie_low_T28Y1;
  wire tie_high_T28Y1;
  wire tie_low_T29Y1;
  wire tie_high_T29Y1;
  wire tie_low_T30Y1;
  wire tie_high_T30Y1;
  wire tie_low_T31Y1;
  wire tie_high_T31Y1;
  wire tie_low_T32Y1;
  wire tie_high_T32Y1;
  wire tie_low_T33Y1;
  wire tie_high_T33Y1;
  wire tie_low_T34Y1;
  wire tie_high_T34Y1;
  wire tie_low_T35Y1;
  wire tie_high_T35Y1;
  wire tie_low_T0Y2;
  wire tie_high_T0Y2;
  wire tie_low_T1Y2;
  wire tie_high_T1Y2;
  wire tie_low_T2Y2;
  wire tie_high_T2Y2;
  wire tie_low_T3Y2;
  wire tie_high_T3Y2;
  wire tie_low_T4Y2;
  wire tie_high_T4Y2;
  wire tie_low_T5Y2;
  wire tie_high_T5Y2;
  wire tie_low_T6Y2;
  wire tie_high_T6Y2;
  wire tie_low_T7Y2;
  wire tie_high_T7Y2;
  wire tie_low_T8Y2;
  wire tie_high_T8Y2;
  wire tie_low_T9Y2;
  wire tie_high_T9Y2;
  wire tie_low_T10Y2;
  wire tie_high_T10Y2;
  wire tie_low_T11Y2;
  wire tie_high_T11Y2;
  wire tie_low_T12Y2;
  wire tie_high_T12Y2;
  wire tie_low_T13Y2;
  wire tie_high_T13Y2;
  wire tie_low_T14Y2;
  wire tie_high_T14Y2;
  wire tie_low_T15Y2;
  wire tie_high_T15Y2;
  wire tie_low_T16Y2;
  wire tie_high_T16Y2;
  wire tie_low_T17Y2;
  wire tie_high_T17Y2;
  wire tie_low_T18Y2;
  wire tie_high_T18Y2;
  wire tie_low_T19Y2;
  wire tie_high_T19Y2;
  wire tie_low_T20Y2;
  wire tie_high_T20Y2;
  wire tie_low_T21Y2;
  wire tie_high_T21Y2;
  wire tie_low_T22Y2;
  wire tie_high_T22Y2;
  wire tie_low_T23Y2;
  wire tie_high_T23Y2;
  wire tie_low_T24Y2;
  wire tie_high_T24Y2;
  wire tie_low_T25Y2;
  wire tie_high_T25Y2;
  wire tie_low_T26Y2;
  wire tie_high_T26Y2;
  wire tie_low_T27Y2;
  wire tie_high_T27Y2;
  wire tie_low_T28Y2;
  wire tie_high_T28Y2;
  wire tie_low_T29Y2;
  wire tie_high_T29Y2;
  wire tie_low_T30Y2;
  wire tie_high_T30Y2;
  wire tie_low_T31Y2;
  wire tie_high_T31Y2;
  wire tie_low_T32Y2;
  wire tie_high_T32Y2;
  wire tie_low_T33Y2;
  wire tie_high_T33Y2;
  wire tie_low_T34Y2;
  wire tie_high_T34Y2;
  wire tie_low_T35Y2;
  wire tie_high_T35Y2;
  wire tie_low_T0Y3;
  wire tie_high_T0Y3;
  wire tie_low_T1Y3;
  wire tie_high_T1Y3;
  wire tie_low_T2Y3;
  wire tie_high_T2Y3;
  wire tie_low_T3Y3;
  wire tie_high_T3Y3;
  wire tie_low_T4Y3;
  wire tie_high_T4Y3;
  wire tie_low_T5Y3;
  wire tie_high_T5Y3;
  wire tie_low_T6Y3;
  wire tie_high_T6Y3;
  wire tie_low_T7Y3;
  wire tie_high_T7Y3;
  wire tie_low_T8Y3;
  wire tie_high_T8Y3;
  wire tie_low_T9Y3;
  wire tie_high_T9Y3;
  wire tie_low_T10Y3;
  wire tie_high_T10Y3;
  wire tie_low_T11Y3;
  wire tie_high_T11Y3;
  wire tie_low_T12Y3;
  wire tie_high_T12Y3;
  wire tie_low_T13Y3;
  wire tie_high_T13Y3;
  wire tie_low_T14Y3;
  wire tie_high_T14Y3;
  wire tie_low_T15Y3;
  wire tie_high_T15Y3;
  wire tie_low_T16Y3;
  wire tie_high_T16Y3;
  wire tie_low_T17Y3;
  wire tie_high_T17Y3;
  wire tie_low_T18Y3;
  wire tie_high_T18Y3;
  wire tie_low_T19Y3;
  wire tie_high_T19Y3;
  wire tie_low_T20Y3;
  wire tie_high_T20Y3;
  wire tie_low_T21Y3;
  wire tie_high_T21Y3;
  wire tie_low_T22Y3;
  wire tie_high_T22Y3;
  wire tie_low_T23Y3;
  wire tie_high_T23Y3;
  wire tie_low_T24Y3;
  wire tie_high_T24Y3;
  wire tie_low_T25Y3;
  wire tie_high_T25Y3;
  wire tie_low_T26Y3;
  wire tie_high_T26Y3;
  wire tie_low_T27Y3;
  wire tie_high_T27Y3;
  wire tie_low_T28Y3;
  wire tie_high_T28Y3;
  wire tie_low_T29Y3;
  wire tie_high_T29Y3;
  wire tie_low_T30Y3;
  wire tie_high_T30Y3;
  wire tie_low_T31Y3;
  wire tie_high_T31Y3;
  wire tie_low_T32Y3;
  wire tie_high_T32Y3;
  wire tie_low_T33Y3;
  wire tie_high_T33Y3;
  wire tie_low_T34Y3;
  wire tie_high_T34Y3;
  wire tie_low_T35Y3;
  wire tie_high_T35Y3;
  wire tie_low_T0Y4;
  wire tie_high_T0Y4;
  wire tie_low_T1Y4;
  wire tie_high_T1Y4;
  wire tie_low_T2Y4;
  wire tie_high_T2Y4;
  wire tie_low_T3Y4;
  wire tie_high_T3Y4;
  wire tie_low_T4Y4;
  wire tie_high_T4Y4;
  wire tie_low_T5Y4;
  wire tie_high_T5Y4;
  wire tie_low_T6Y4;
  wire tie_high_T6Y4;
  wire tie_low_T7Y4;
  wire tie_high_T7Y4;
  wire tie_low_T8Y4;
  wire tie_high_T8Y4;
  wire tie_low_T9Y4;
  wire tie_high_T9Y4;
  wire tie_low_T10Y4;
  wire tie_high_T10Y4;
  wire tie_low_T11Y4;
  wire tie_high_T11Y4;
  wire tie_low_T12Y4;
  wire tie_high_T12Y4;
  wire tie_low_T13Y4;
  wire tie_high_T13Y4;
  wire tie_low_T14Y4;
  wire tie_high_T14Y4;
  wire tie_low_T15Y4;
  wire tie_high_T15Y4;
  wire tie_low_T16Y4;
  wire tie_high_T16Y4;
  wire tie_low_T17Y4;
  wire tie_high_T17Y4;
  wire tie_low_T18Y4;
  wire tie_high_T18Y4;
  wire tie_low_T19Y4;
  wire tie_high_T19Y4;
  wire tie_low_T20Y4;
  wire tie_high_T20Y4;
  wire tie_low_T21Y4;
  wire tie_high_T21Y4;
  wire tie_low_T22Y4;
  wire tie_high_T22Y4;
  wire tie_low_T23Y4;
  wire tie_high_T23Y4;
  wire tie_low_T24Y4;
  wire tie_high_T24Y4;
  wire tie_low_T25Y4;
  wire tie_high_T25Y4;
  wire tie_low_T26Y4;
  wire tie_high_T26Y4;
  wire tie_low_T27Y4;
  wire tie_high_T27Y4;
  wire tie_low_T28Y4;
  wire tie_high_T28Y4;
  wire tie_low_T29Y4;
  wire tie_high_T29Y4;
  wire tie_low_T30Y4;
  wire tie_high_T30Y4;
  wire tie_low_T31Y4;
  wire tie_high_T31Y4;
  wire tie_low_T32Y4;
  wire tie_high_T32Y4;
  wire tie_low_T33Y4;
  wire tie_high_T33Y4;
  wire tie_low_T34Y4;
  wire tie_high_T34Y4;
  wire tie_low_T35Y4;
  wire tie_high_T35Y4;
  wire tie_low_T0Y5;
  wire tie_high_T0Y5;
  wire tie_low_T1Y5;
  wire tie_high_T1Y5;
  wire tie_low_T2Y5;
  wire tie_high_T2Y5;
  wire tie_low_T3Y5;
  wire tie_high_T3Y5;
  wire tie_low_T4Y5;
  wire tie_high_T4Y5;
  wire tie_low_T5Y5;
  wire tie_high_T5Y5;
  wire tie_low_T6Y5;
  wire tie_high_T6Y5;
  wire tie_low_T7Y5;
  wire tie_high_T7Y5;
  wire tie_low_T8Y5;
  wire tie_high_T8Y5;
  wire tie_low_T9Y5;
  wire tie_high_T9Y5;
  wire tie_low_T10Y5;
  wire tie_high_T10Y5;
  wire tie_low_T11Y5;
  wire tie_high_T11Y5;
  wire tie_low_T12Y5;
  wire tie_high_T12Y5;
  wire tie_low_T13Y5;
  wire tie_high_T13Y5;
  wire tie_low_T14Y5;
  wire tie_high_T14Y5;
  wire tie_low_T15Y5;
  wire tie_high_T15Y5;
  wire tie_low_T16Y5;
  wire tie_high_T16Y5;
  wire tie_low_T17Y5;
  wire tie_high_T17Y5;
  wire tie_low_T18Y5;
  wire tie_high_T18Y5;
  wire tie_low_T19Y5;
  wire tie_high_T19Y5;
  wire tie_low_T20Y5;
  wire tie_high_T20Y5;
  wire tie_low_T21Y5;
  wire tie_high_T21Y5;
  wire tie_low_T22Y5;
  wire tie_high_T22Y5;
  wire tie_low_T23Y5;
  wire tie_high_T23Y5;
  wire tie_low_T24Y5;
  wire tie_high_T24Y5;
  wire tie_low_T25Y5;
  wire tie_high_T25Y5;
  wire tie_low_T26Y5;
  wire tie_high_T26Y5;
  wire tie_low_T27Y5;
  wire tie_high_T27Y5;
  wire tie_low_T28Y5;
  wire tie_high_T28Y5;
  wire tie_low_T29Y5;
  wire tie_high_T29Y5;
  wire tie_low_T30Y5;
  wire tie_high_T30Y5;
  wire tie_low_T31Y5;
  wire tie_high_T31Y5;
  wire tie_low_T32Y5;
  wire tie_high_T32Y5;
  wire tie_low_T33Y5;
  wire tie_high_T33Y5;
  wire tie_low_T34Y5;
  wire tie_high_T34Y5;
  wire tie_low_T35Y5;
  wire tie_high_T35Y5;
  wire tie_low_T0Y6;
  wire tie_high_T0Y6;
  wire tie_low_T1Y6;
  wire tie_high_T1Y6;
  wire tie_low_T2Y6;
  wire tie_high_T2Y6;
  wire tie_low_T3Y6;
  wire tie_high_T3Y6;
  wire tie_low_T4Y6;
  wire tie_high_T4Y6;
  wire tie_low_T5Y6;
  wire tie_high_T5Y6;
  wire tie_low_T6Y6;
  wire tie_high_T6Y6;
  wire tie_low_T7Y6;
  wire tie_high_T7Y6;
  wire tie_low_T8Y6;
  wire tie_high_T8Y6;
  wire tie_low_T9Y6;
  wire tie_high_T9Y6;
  wire tie_low_T10Y6;
  wire tie_high_T10Y6;
  wire tie_low_T11Y6;
  wire tie_high_T11Y6;
  wire tie_low_T12Y6;
  wire tie_high_T12Y6;
  wire tie_low_T13Y6;
  wire tie_high_T13Y6;
  wire tie_low_T14Y6;
  wire tie_high_T14Y6;
  wire tie_low_T15Y6;
  wire tie_high_T15Y6;
  wire tie_low_T16Y6;
  wire tie_high_T16Y6;
  wire tie_low_T17Y6;
  wire tie_high_T17Y6;
  wire tie_low_T18Y6;
  wire tie_high_T18Y6;
  wire tie_low_T19Y6;
  wire tie_high_T19Y6;
  wire tie_low_T20Y6;
  wire tie_high_T20Y6;
  wire tie_low_T21Y6;
  wire tie_high_T21Y6;
  wire tie_low_T22Y6;
  wire tie_high_T22Y6;
  wire tie_low_T23Y6;
  wire tie_high_T23Y6;
  wire tie_low_T24Y6;
  wire tie_high_T24Y6;
  wire tie_low_T25Y6;
  wire tie_high_T25Y6;
  wire tie_low_T26Y6;
  wire tie_high_T26Y6;
  wire tie_low_T27Y6;
  wire tie_high_T27Y6;
  wire tie_low_T28Y6;
  wire tie_high_T28Y6;
  wire tie_low_T29Y6;
  wire tie_high_T29Y6;
  wire tie_low_T30Y6;
  wire tie_high_T30Y6;
  wire tie_low_T31Y6;
  wire tie_high_T31Y6;
  wire tie_low_T32Y6;
  wire tie_high_T32Y6;
  wire tie_low_T33Y6;
  wire tie_high_T33Y6;
  wire tie_low_T34Y6;
  wire tie_high_T34Y6;
  wire tie_low_T35Y6;
  wire tie_high_T35Y6;
  wire tie_low_T0Y7;
  wire tie_high_T0Y7;
  wire tie_low_T1Y7;
  wire tie_high_T1Y7;
  wire tie_low_T2Y7;
  wire tie_high_T2Y7;
  wire tie_low_T3Y7;
  wire tie_high_T3Y7;
  wire tie_low_T4Y7;
  wire tie_high_T4Y7;
  wire tie_low_T5Y7;
  wire tie_high_T5Y7;
  wire tie_low_T6Y7;
  wire tie_high_T6Y7;
  wire tie_low_T7Y7;
  wire tie_high_T7Y7;
  wire tie_low_T8Y7;
  wire tie_high_T8Y7;
  wire tie_low_T9Y7;
  wire tie_high_T9Y7;
  wire tie_low_T10Y7;
  wire tie_high_T10Y7;
  wire tie_low_T11Y7;
  wire tie_high_T11Y7;
  wire tie_low_T12Y7;
  wire tie_high_T12Y7;
  wire tie_low_T13Y7;
  wire tie_high_T13Y7;
  wire tie_low_T14Y7;
  wire tie_high_T14Y7;
  wire tie_low_T15Y7;
  wire tie_high_T15Y7;
  wire tie_low_T16Y7;
  wire tie_high_T16Y7;
  wire tie_low_T17Y7;
  wire tie_high_T17Y7;
  wire tie_low_T18Y7;
  wire tie_high_T18Y7;
  wire tie_low_T19Y7;
  wire tie_high_T19Y7;
  wire tie_low_T20Y7;
  wire tie_high_T20Y7;
  wire tie_low_T21Y7;
  wire tie_high_T21Y7;
  wire tie_low_T22Y7;
  wire tie_high_T22Y7;
  wire tie_low_T23Y7;
  wire tie_high_T23Y7;
  wire tie_low_T24Y7;
  wire tie_high_T24Y7;
  wire tie_low_T25Y7;
  wire tie_high_T25Y7;
  wire tie_low_T26Y7;
  wire tie_high_T26Y7;
  wire tie_low_T27Y7;
  wire tie_high_T27Y7;
  wire tie_low_T28Y7;
  wire tie_high_T28Y7;
  wire tie_low_T29Y7;
  wire tie_high_T29Y7;
  wire tie_low_T30Y7;
  wire tie_high_T30Y7;
  wire tie_low_T31Y7;
  wire tie_high_T31Y7;
  wire tie_low_T32Y7;
  wire tie_high_T32Y7;
  wire tie_low_T33Y7;
  wire tie_high_T33Y7;
  wire tie_low_T34Y7;
  wire tie_high_T34Y7;
  wire tie_low_T35Y7;
  wire tie_high_T35Y7;
  wire tie_low_T0Y8;
  wire tie_high_T0Y8;
  wire tie_low_T1Y8;
  wire tie_high_T1Y8;
  wire tie_low_T2Y8;
  wire tie_high_T2Y8;
  wire tie_low_T3Y8;
  wire tie_high_T3Y8;
  wire tie_low_T4Y8;
  wire tie_high_T4Y8;
  wire tie_low_T5Y8;
  wire tie_high_T5Y8;
  wire tie_low_T6Y8;
  wire tie_high_T6Y8;
  wire tie_low_T7Y8;
  wire tie_high_T7Y8;
  wire tie_low_T8Y8;
  wire tie_high_T8Y8;
  wire tie_low_T9Y8;
  wire tie_high_T9Y8;
  wire tie_low_T10Y8;
  wire tie_high_T10Y8;
  wire tie_low_T11Y8;
  wire tie_high_T11Y8;
  wire tie_low_T12Y8;
  wire tie_high_T12Y8;
  wire tie_low_T13Y8;
  wire tie_high_T13Y8;
  wire tie_low_T14Y8;
  wire tie_high_T14Y8;
  wire tie_low_T15Y8;
  wire tie_high_T15Y8;
  wire tie_low_T16Y8;
  wire tie_high_T16Y8;
  wire tie_low_T17Y8;
  wire tie_high_T17Y8;
  wire tie_low_T18Y8;
  wire tie_high_T18Y8;
  wire tie_low_T19Y8;
  wire tie_high_T19Y8;
  wire tie_low_T20Y8;
  wire tie_high_T20Y8;
  wire tie_low_T21Y8;
  wire tie_high_T21Y8;
  wire tie_low_T22Y8;
  wire tie_high_T22Y8;
  wire tie_low_T23Y8;
  wire tie_high_T23Y8;
  wire tie_low_T24Y8;
  wire tie_high_T24Y8;
  wire tie_low_T25Y8;
  wire tie_high_T25Y8;
  wire tie_low_T26Y8;
  wire tie_high_T26Y8;
  wire tie_low_T27Y8;
  wire tie_high_T27Y8;
  wire tie_low_T28Y8;
  wire tie_high_T28Y8;
  wire tie_low_T29Y8;
  wire tie_high_T29Y8;
  wire tie_low_T30Y8;
  wire tie_high_T30Y8;
  wire tie_low_T31Y8;
  wire tie_high_T31Y8;
  wire tie_low_T32Y8;
  wire tie_high_T32Y8;
  wire tie_low_T33Y8;
  wire tie_high_T33Y8;
  wire tie_low_T34Y8;
  wire tie_high_T34Y8;
  wire tie_low_T35Y8;
  wire tie_high_T35Y8;
  wire tie_low_T0Y9;
  wire tie_high_T0Y9;
  wire tie_low_T1Y9;
  wire tie_high_T1Y9;
  wire tie_low_T2Y9;
  wire tie_high_T2Y9;
  wire tie_low_T3Y9;
  wire tie_high_T3Y9;
  wire tie_low_T4Y9;
  wire tie_high_T4Y9;
  wire tie_low_T5Y9;
  wire tie_high_T5Y9;
  wire tie_low_T6Y9;
  wire tie_high_T6Y9;
  wire tie_low_T7Y9;
  wire tie_high_T7Y9;
  wire tie_low_T8Y9;
  wire tie_high_T8Y9;
  wire tie_low_T9Y9;
  wire tie_high_T9Y9;
  wire tie_low_T10Y9;
  wire tie_high_T10Y9;
  wire tie_low_T11Y9;
  wire tie_high_T11Y9;
  wire tie_low_T12Y9;
  wire tie_high_T12Y9;
  wire tie_low_T13Y9;
  wire tie_high_T13Y9;
  wire tie_low_T14Y9;
  wire tie_high_T14Y9;
  wire tie_low_T15Y9;
  wire tie_high_T15Y9;
  wire tie_low_T16Y9;
  wire tie_high_T16Y9;
  wire tie_low_T17Y9;
  wire tie_high_T17Y9;
  wire tie_low_T18Y9;
  wire tie_high_T18Y9;
  wire tie_low_T19Y9;
  wire tie_high_T19Y9;
  wire tie_low_T20Y9;
  wire tie_high_T20Y9;
  wire tie_low_T21Y9;
  wire tie_high_T21Y9;
  wire tie_low_T22Y9;
  wire tie_high_T22Y9;
  wire tie_low_T23Y9;
  wire tie_high_T23Y9;
  wire tie_low_T24Y9;
  wire tie_high_T24Y9;
  wire tie_low_T25Y9;
  wire tie_high_T25Y9;
  wire tie_low_T26Y9;
  wire tie_high_T26Y9;
  wire tie_low_T27Y9;
  wire tie_high_T27Y9;
  wire tie_low_T28Y9;
  wire tie_high_T28Y9;
  wire tie_low_T29Y9;
  wire tie_high_T29Y9;
  wire tie_low_T30Y9;
  wire tie_high_T30Y9;
  wire tie_low_T31Y9;
  wire tie_high_T31Y9;
  wire tie_low_T32Y9;
  wire tie_high_T32Y9;
  wire tie_low_T33Y9;
  wire tie_high_T33Y9;
  wire tie_low_T34Y9;
  wire tie_high_T34Y9;
  wire tie_low_T35Y9;
  wire tie_high_T35Y9;
  wire tie_low_T0Y10;
  wire tie_high_T0Y10;
  wire tie_low_T1Y10;
  wire tie_high_T1Y10;
  wire tie_low_T2Y10;
  wire tie_high_T2Y10;
  wire tie_low_T3Y10;
  wire tie_high_T3Y10;
  wire tie_low_T4Y10;
  wire tie_high_T4Y10;
  wire tie_low_T5Y10;
  wire tie_high_T5Y10;
  wire tie_low_T6Y10;
  wire tie_high_T6Y10;
  wire tie_low_T7Y10;
  wire tie_high_T7Y10;
  wire tie_low_T8Y10;
  wire tie_high_T8Y10;
  wire tie_low_T9Y10;
  wire tie_high_T9Y10;
  wire tie_low_T10Y10;
  wire tie_high_T10Y10;
  wire tie_low_T11Y10;
  wire tie_high_T11Y10;
  wire tie_low_T12Y10;
  wire tie_high_T12Y10;
  wire tie_low_T13Y10;
  wire tie_high_T13Y10;
  wire tie_low_T14Y10;
  wire tie_high_T14Y10;
  wire tie_low_T15Y10;
  wire tie_high_T15Y10;
  wire tie_low_T16Y10;
  wire tie_high_T16Y10;
  wire tie_low_T17Y10;
  wire tie_high_T17Y10;
  wire tie_low_T18Y10;
  wire tie_high_T18Y10;
  wire tie_low_T19Y10;
  wire tie_high_T19Y10;
  wire tie_low_T20Y10;
  wire tie_high_T20Y10;
  wire tie_low_T21Y10;
  wire tie_high_T21Y10;
  wire tie_low_T22Y10;
  wire tie_high_T22Y10;
  wire tie_low_T23Y10;
  wire tie_high_T23Y10;
  wire tie_low_T24Y10;
  wire tie_high_T24Y10;
  wire tie_low_T25Y10;
  wire tie_high_T25Y10;
  wire tie_low_T26Y10;
  wire tie_high_T26Y10;
  wire tie_low_T27Y10;
  wire tie_high_T27Y10;
  wire tie_low_T28Y10;
  wire tie_high_T28Y10;
  wire tie_low_T29Y10;
  wire tie_high_T29Y10;
  wire tie_low_T30Y10;
  wire tie_high_T30Y10;
  wire tie_low_T31Y10;
  wire tie_high_T31Y10;
  wire tie_low_T32Y10;
  wire tie_high_T32Y10;
  wire tie_low_T33Y10;
  wire tie_high_T33Y10;
  wire tie_low_T34Y10;
  wire tie_high_T34Y10;
  wire tie_low_T35Y10;
  wire tie_high_T35Y10;
  wire tie_low_T0Y11;
  wire tie_high_T0Y11;
  wire tie_low_T1Y11;
  wire tie_high_T1Y11;
  wire tie_low_T2Y11;
  wire tie_high_T2Y11;
  wire tie_low_T3Y11;
  wire tie_high_T3Y11;
  wire tie_low_T4Y11;
  wire tie_high_T4Y11;
  wire tie_low_T5Y11;
  wire tie_high_T5Y11;
  wire tie_low_T6Y11;
  wire tie_high_T6Y11;
  wire tie_low_T7Y11;
  wire tie_high_T7Y11;
  wire tie_low_T8Y11;
  wire tie_high_T8Y11;
  wire tie_low_T9Y11;
  wire tie_high_T9Y11;
  wire tie_low_T10Y11;
  wire tie_high_T10Y11;
  wire tie_low_T11Y11;
  wire tie_high_T11Y11;
  wire tie_low_T12Y11;
  wire tie_high_T12Y11;
  wire tie_low_T13Y11;
  wire tie_high_T13Y11;
  wire tie_low_T14Y11;
  wire tie_high_T14Y11;
  wire tie_low_T15Y11;
  wire tie_high_T15Y11;
  wire tie_low_T16Y11;
  wire tie_high_T16Y11;
  wire tie_low_T17Y11;
  wire tie_high_T17Y11;
  wire tie_low_T18Y11;
  wire tie_high_T18Y11;
  wire tie_low_T19Y11;
  wire tie_high_T19Y11;
  wire tie_low_T20Y11;
  wire tie_high_T20Y11;
  wire tie_low_T21Y11;
  wire tie_high_T21Y11;
  wire tie_low_T22Y11;
  wire tie_high_T22Y11;
  wire tie_low_T23Y11;
  wire tie_high_T23Y11;
  wire tie_low_T24Y11;
  wire tie_high_T24Y11;
  wire tie_low_T25Y11;
  wire tie_high_T25Y11;
  wire tie_low_T26Y11;
  wire tie_high_T26Y11;
  wire tie_low_T27Y11;
  wire tie_high_T27Y11;
  wire tie_low_T28Y11;
  wire tie_high_T28Y11;
  wire tie_low_T29Y11;
  wire tie_high_T29Y11;
  wire tie_low_T30Y11;
  wire tie_high_T30Y11;
  wire tie_low_T31Y11;
  wire tie_high_T31Y11;
  wire tie_low_T32Y11;
  wire tie_high_T32Y11;
  wire tie_low_T33Y11;
  wire tie_high_T33Y11;
  wire tie_low_T34Y11;
  wire tie_high_T34Y11;
  wire tie_low_T35Y11;
  wire tie_high_T35Y11;
  wire tie_low_T0Y12;
  wire tie_high_T0Y12;
  wire tie_low_T1Y12;
  wire tie_high_T1Y12;
  wire tie_low_T2Y12;
  wire tie_high_T2Y12;
  wire tie_low_T3Y12;
  wire tie_high_T3Y12;
  wire tie_low_T4Y12;
  wire tie_high_T4Y12;
  wire tie_low_T5Y12;
  wire tie_high_T5Y12;
  wire tie_low_T6Y12;
  wire tie_high_T6Y12;
  wire tie_low_T7Y12;
  wire tie_high_T7Y12;
  wire tie_low_T8Y12;
  wire tie_high_T8Y12;
  wire tie_low_T9Y12;
  wire tie_high_T9Y12;
  wire tie_low_T10Y12;
  wire tie_high_T10Y12;
  wire tie_low_T11Y12;
  wire tie_high_T11Y12;
  wire tie_low_T12Y12;
  wire tie_high_T12Y12;
  wire tie_low_T13Y12;
  wire tie_high_T13Y12;
  wire tie_low_T14Y12;
  wire tie_high_T14Y12;
  wire tie_low_T15Y12;
  wire tie_high_T15Y12;
  wire tie_low_T16Y12;
  wire tie_high_T16Y12;
  wire tie_low_T17Y12;
  wire tie_high_T17Y12;
  wire tie_low_T18Y12;
  wire tie_high_T18Y12;
  wire tie_low_T19Y12;
  wire tie_high_T19Y12;
  wire tie_low_T20Y12;
  wire tie_high_T20Y12;
  wire tie_low_T21Y12;
  wire tie_high_T21Y12;
  wire tie_low_T22Y12;
  wire tie_high_T22Y12;
  wire tie_low_T23Y12;
  wire tie_high_T23Y12;
  wire tie_low_T24Y12;
  wire tie_high_T24Y12;
  wire tie_low_T25Y12;
  wire tie_high_T25Y12;
  wire tie_low_T26Y12;
  wire tie_high_T26Y12;
  wire tie_low_T27Y12;
  wire tie_high_T27Y12;
  wire tie_low_T28Y12;
  wire tie_high_T28Y12;
  wire tie_low_T29Y12;
  wire tie_high_T29Y12;
  wire tie_low_T30Y12;
  wire tie_high_T30Y12;
  wire tie_low_T31Y12;
  wire tie_high_T31Y12;
  wire tie_low_T32Y12;
  wire tie_high_T32Y12;
  wire tie_low_T33Y12;
  wire tie_high_T33Y12;
  wire tie_low_T34Y12;
  wire tie_high_T34Y12;
  wire tie_low_T35Y12;
  wire tie_high_T35Y12;
  wire tie_low_T0Y13;
  wire tie_high_T0Y13;
  wire tie_low_T1Y13;
  wire tie_high_T1Y13;
  wire tie_low_T2Y13;
  wire tie_high_T2Y13;
  wire tie_low_T3Y13;
  wire tie_high_T3Y13;
  wire tie_low_T4Y13;
  wire tie_high_T4Y13;
  wire tie_low_T5Y13;
  wire tie_high_T5Y13;
  wire tie_low_T6Y13;
  wire tie_high_T6Y13;
  wire tie_low_T7Y13;
  wire tie_high_T7Y13;
  wire tie_low_T8Y13;
  wire tie_high_T8Y13;
  wire tie_low_T9Y13;
  wire tie_high_T9Y13;
  wire tie_low_T10Y13;
  wire tie_high_T10Y13;
  wire tie_low_T11Y13;
  wire tie_high_T11Y13;
  wire tie_low_T12Y13;
  wire tie_high_T12Y13;
  wire tie_low_T13Y13;
  wire tie_high_T13Y13;
  wire tie_low_T14Y13;
  wire tie_high_T14Y13;
  wire tie_low_T15Y13;
  wire tie_high_T15Y13;
  wire tie_low_T16Y13;
  wire tie_high_T16Y13;
  wire tie_low_T17Y13;
  wire tie_high_T17Y13;
  wire tie_low_T18Y13;
  wire tie_high_T18Y13;
  wire tie_low_T19Y13;
  wire tie_high_T19Y13;
  wire tie_low_T20Y13;
  wire tie_high_T20Y13;
  wire tie_low_T21Y13;
  wire tie_high_T21Y13;
  wire tie_low_T22Y13;
  wire tie_high_T22Y13;
  wire tie_low_T23Y13;
  wire tie_high_T23Y13;
  wire tie_low_T24Y13;
  wire tie_high_T24Y13;
  wire tie_low_T25Y13;
  wire tie_high_T25Y13;
  wire tie_low_T26Y13;
  wire tie_high_T26Y13;
  wire tie_low_T27Y13;
  wire tie_high_T27Y13;
  wire tie_low_T28Y13;
  wire tie_high_T28Y13;
  wire tie_low_T29Y13;
  wire tie_high_T29Y13;
  wire tie_low_T30Y13;
  wire tie_high_T30Y13;
  wire tie_low_T31Y13;
  wire tie_high_T31Y13;
  wire tie_low_T32Y13;
  wire tie_high_T32Y13;
  wire tie_low_T33Y13;
  wire tie_high_T33Y13;
  wire tie_low_T34Y13;
  wire tie_high_T34Y13;
  wire tie_low_T35Y13;
  wire tie_high_T35Y13;
  wire tie_low_T0Y14;
  wire tie_high_T0Y14;
  wire tie_low_T1Y14;
  wire tie_high_T1Y14;
  wire tie_low_T2Y14;
  wire tie_high_T2Y14;
  wire tie_low_T3Y14;
  wire tie_high_T3Y14;
  wire tie_low_T4Y14;
  wire tie_high_T4Y14;
  wire tie_low_T5Y14;
  wire tie_high_T5Y14;
  wire tie_low_T6Y14;
  wire tie_high_T6Y14;
  wire tie_low_T7Y14;
  wire tie_high_T7Y14;
  wire tie_low_T8Y14;
  wire tie_high_T8Y14;
  wire tie_low_T9Y14;
  wire tie_high_T9Y14;
  wire tie_low_T10Y14;
  wire tie_high_T10Y14;
  wire tie_low_T11Y14;
  wire tie_high_T11Y14;
  wire tie_low_T12Y14;
  wire tie_high_T12Y14;
  wire tie_low_T13Y14;
  wire tie_high_T13Y14;
  wire tie_low_T14Y14;
  wire tie_high_T14Y14;
  wire tie_low_T15Y14;
  wire tie_high_T15Y14;
  wire tie_low_T16Y14;
  wire tie_high_T16Y14;
  wire tie_low_T17Y14;
  wire tie_high_T17Y14;
  wire tie_low_T18Y14;
  wire tie_high_T18Y14;
  wire tie_low_T19Y14;
  wire tie_high_T19Y14;
  wire tie_low_T20Y14;
  wire tie_high_T20Y14;
  wire tie_low_T21Y14;
  wire tie_high_T21Y14;
  wire tie_low_T22Y14;
  wire tie_high_T22Y14;
  wire tie_low_T23Y14;
  wire tie_high_T23Y14;
  wire tie_low_T24Y14;
  wire tie_high_T24Y14;
  wire tie_low_T25Y14;
  wire tie_high_T25Y14;
  wire tie_low_T26Y14;
  wire tie_high_T26Y14;
  wire tie_low_T27Y14;
  wire tie_high_T27Y14;
  wire tie_low_T28Y14;
  wire tie_high_T28Y14;
  wire tie_low_T29Y14;
  wire tie_high_T29Y14;
  wire tie_low_T30Y14;
  wire tie_high_T30Y14;
  wire tie_low_T31Y14;
  wire tie_high_T31Y14;
  wire tie_low_T32Y14;
  wire tie_high_T32Y14;
  wire tie_low_T33Y14;
  wire tie_high_T33Y14;
  wire tie_low_T34Y14;
  wire tie_high_T34Y14;
  wire tie_low_T35Y14;
  wire tie_high_T35Y14;
  wire tie_low_T0Y15;
  wire tie_high_T0Y15;
  wire tie_low_T1Y15;
  wire tie_high_T1Y15;
  wire tie_low_T2Y15;
  wire tie_high_T2Y15;
  wire tie_low_T3Y15;
  wire tie_high_T3Y15;
  wire tie_low_T4Y15;
  wire tie_high_T4Y15;
  wire tie_low_T5Y15;
  wire tie_high_T5Y15;
  wire tie_low_T6Y15;
  wire tie_high_T6Y15;
  wire tie_low_T7Y15;
  wire tie_high_T7Y15;
  wire tie_low_T8Y15;
  wire tie_high_T8Y15;
  wire tie_low_T9Y15;
  wire tie_high_T9Y15;
  wire tie_low_T10Y15;
  wire tie_high_T10Y15;
  wire tie_low_T11Y15;
  wire tie_high_T11Y15;
  wire tie_low_T12Y15;
  wire tie_high_T12Y15;
  wire tie_low_T13Y15;
  wire tie_high_T13Y15;
  wire tie_low_T14Y15;
  wire tie_high_T14Y15;
  wire tie_low_T15Y15;
  wire tie_high_T15Y15;
  wire tie_low_T16Y15;
  wire tie_high_T16Y15;
  wire tie_low_T17Y15;
  wire tie_high_T17Y15;
  wire tie_low_T18Y15;
  wire tie_high_T18Y15;
  wire tie_low_T19Y15;
  wire tie_high_T19Y15;
  wire tie_low_T20Y15;
  wire tie_high_T20Y15;
  wire tie_low_T21Y15;
  wire tie_high_T21Y15;
  wire tie_low_T22Y15;
  wire tie_high_T22Y15;
  wire tie_low_T23Y15;
  wire tie_high_T23Y15;
  wire tie_low_T24Y15;
  wire tie_high_T24Y15;
  wire tie_low_T25Y15;
  wire tie_high_T25Y15;
  wire tie_low_T26Y15;
  wire tie_high_T26Y15;
  wire tie_low_T27Y15;
  wire tie_high_T27Y15;
  wire tie_low_T28Y15;
  wire tie_high_T28Y15;
  wire tie_low_T29Y15;
  wire tie_high_T29Y15;
  wire tie_low_T30Y15;
  wire tie_high_T30Y15;
  wire tie_low_T31Y15;
  wire tie_high_T31Y15;
  wire tie_low_T32Y15;
  wire tie_high_T32Y15;
  wire tie_low_T33Y15;
  wire tie_high_T33Y15;
  wire tie_low_T34Y15;
  wire tie_high_T34Y15;
  wire tie_low_T35Y15;
  wire tie_high_T35Y15;
  wire tie_low_T0Y16;
  wire tie_high_T0Y16;
  wire tie_low_T1Y16;
  wire tie_high_T1Y16;
  wire tie_low_T2Y16;
  wire tie_high_T2Y16;
  wire tie_low_T3Y16;
  wire tie_high_T3Y16;
  wire tie_low_T4Y16;
  wire tie_high_T4Y16;
  wire tie_low_T5Y16;
  wire tie_high_T5Y16;
  wire tie_low_T6Y16;
  wire tie_high_T6Y16;
  wire tie_low_T7Y16;
  wire tie_high_T7Y16;
  wire tie_low_T8Y16;
  wire tie_high_T8Y16;
  wire tie_low_T9Y16;
  wire tie_high_T9Y16;
  wire tie_low_T10Y16;
  wire tie_high_T10Y16;
  wire tie_low_T11Y16;
  wire tie_high_T11Y16;
  wire tie_low_T12Y16;
  wire tie_high_T12Y16;
  wire tie_low_T13Y16;
  wire tie_high_T13Y16;
  wire tie_low_T14Y16;
  wire tie_high_T14Y16;
  wire tie_low_T15Y16;
  wire tie_high_T15Y16;
  wire tie_low_T16Y16;
  wire tie_high_T16Y16;
  wire tie_low_T17Y16;
  wire tie_high_T17Y16;
  wire tie_low_T18Y16;
  wire tie_high_T18Y16;
  wire tie_low_T19Y16;
  wire tie_high_T19Y16;
  wire tie_low_T20Y16;
  wire tie_high_T20Y16;
  wire tie_low_T21Y16;
  wire tie_high_T21Y16;
  wire tie_low_T22Y16;
  wire tie_high_T22Y16;
  wire tie_low_T23Y16;
  wire tie_high_T23Y16;
  wire tie_low_T24Y16;
  wire tie_high_T24Y16;
  wire tie_low_T25Y16;
  wire tie_high_T25Y16;
  wire tie_low_T26Y16;
  wire tie_high_T26Y16;
  wire tie_low_T27Y16;
  wire tie_high_T27Y16;
  wire tie_low_T28Y16;
  wire tie_high_T28Y16;
  wire tie_low_T29Y16;
  wire tie_high_T29Y16;
  wire tie_low_T30Y16;
  wire tie_high_T30Y16;
  wire tie_low_T31Y16;
  wire tie_high_T31Y16;
  wire tie_low_T32Y16;
  wire tie_high_T32Y16;
  wire tie_low_T33Y16;
  wire tie_high_T33Y16;
  wire tie_low_T34Y16;
  wire tie_high_T34Y16;
  wire tie_low_T35Y16;
  wire tie_high_T35Y16;
  wire tie_low_T0Y17;
  wire tie_high_T0Y17;
  wire tie_low_T1Y17;
  wire tie_high_T1Y17;
  wire tie_low_T2Y17;
  wire tie_high_T2Y17;
  wire tie_low_T3Y17;
  wire tie_high_T3Y17;
  wire tie_low_T4Y17;
  wire tie_high_T4Y17;
  wire tie_low_T5Y17;
  wire tie_high_T5Y17;
  wire tie_low_T6Y17;
  wire tie_high_T6Y17;
  wire tie_low_T7Y17;
  wire tie_high_T7Y17;
  wire tie_low_T8Y17;
  wire tie_high_T8Y17;
  wire tie_low_T9Y17;
  wire tie_high_T9Y17;
  wire tie_low_T10Y17;
  wire tie_high_T10Y17;
  wire tie_low_T11Y17;
  wire tie_high_T11Y17;
  wire tie_low_T12Y17;
  wire tie_high_T12Y17;
  wire tie_low_T13Y17;
  wire tie_high_T13Y17;
  wire tie_low_T14Y17;
  wire tie_high_T14Y17;
  wire tie_low_T15Y17;
  wire tie_high_T15Y17;
  wire tie_low_T16Y17;
  wire tie_high_T16Y17;
  wire tie_low_T17Y17;
  wire tie_high_T17Y17;
  wire tie_low_T18Y17;
  wire tie_high_T18Y17;
  wire tie_low_T19Y17;
  wire tie_high_T19Y17;
  wire tie_low_T20Y17;
  wire tie_high_T20Y17;
  wire tie_low_T21Y17;
  wire tie_high_T21Y17;
  wire tie_low_T22Y17;
  wire tie_high_T22Y17;
  wire tie_low_T23Y17;
  wire tie_high_T23Y17;
  wire tie_low_T24Y17;
  wire tie_high_T24Y17;
  wire tie_low_T25Y17;
  wire tie_high_T25Y17;
  wire tie_low_T26Y17;
  wire tie_high_T26Y17;
  wire tie_low_T27Y17;
  wire tie_high_T27Y17;
  wire tie_low_T28Y17;
  wire tie_high_T28Y17;
  wire tie_low_T29Y17;
  wire tie_high_T29Y17;
  wire tie_low_T30Y17;
  wire tie_high_T30Y17;
  wire tie_low_T31Y17;
  wire tie_high_T31Y17;
  wire tie_low_T32Y17;
  wire tie_high_T32Y17;
  wire tie_low_T33Y17;
  wire tie_high_T33Y17;
  wire tie_low_T34Y17;
  wire tie_high_T34Y17;
  wire tie_low_T35Y17;
  wire tie_high_T35Y17;
  wire tie_low_T0Y18;
  wire tie_high_T0Y18;
  wire tie_low_T1Y18;
  wire tie_high_T1Y18;
  wire tie_low_T2Y18;
  wire tie_high_T2Y18;
  wire tie_low_T3Y18;
  wire tie_high_T3Y18;
  wire tie_low_T4Y18;
  wire tie_high_T4Y18;
  wire tie_low_T5Y18;
  wire tie_high_T5Y18;
  wire tie_low_T6Y18;
  wire tie_high_T6Y18;
  wire tie_low_T7Y18;
  wire tie_high_T7Y18;
  wire tie_low_T8Y18;
  wire tie_high_T8Y18;
  wire tie_low_T9Y18;
  wire tie_high_T9Y18;
  wire tie_low_T10Y18;
  wire tie_high_T10Y18;
  wire tie_low_T11Y18;
  wire tie_high_T11Y18;
  wire tie_low_T12Y18;
  wire tie_high_T12Y18;
  wire tie_low_T13Y18;
  wire tie_high_T13Y18;
  wire tie_low_T14Y18;
  wire tie_high_T14Y18;
  wire tie_low_T15Y18;
  wire tie_high_T15Y18;
  wire tie_low_T16Y18;
  wire tie_high_T16Y18;
  wire tie_low_T17Y18;
  wire tie_high_T17Y18;
  wire tie_low_T18Y18;
  wire tie_high_T18Y18;
  wire tie_low_T19Y18;
  wire tie_high_T19Y18;
  wire tie_low_T20Y18;
  wire tie_high_T20Y18;
  wire tie_low_T21Y18;
  wire tie_high_T21Y18;
  wire tie_low_T22Y18;
  wire tie_high_T22Y18;
  wire tie_low_T23Y18;
  wire tie_high_T23Y18;
  wire tie_low_T24Y18;
  wire tie_high_T24Y18;
  wire tie_low_T25Y18;
  wire tie_high_T25Y18;
  wire tie_low_T26Y18;
  wire tie_high_T26Y18;
  wire tie_low_T27Y18;
  wire tie_high_T27Y18;
  wire tie_low_T28Y18;
  wire tie_high_T28Y18;
  wire tie_low_T29Y18;
  wire tie_high_T29Y18;
  wire tie_low_T30Y18;
  wire tie_high_T30Y18;
  wire tie_low_T31Y18;
  wire tie_high_T31Y18;
  wire tie_low_T32Y18;
  wire tie_high_T32Y18;
  wire tie_low_T33Y18;
  wire tie_high_T33Y18;
  wire tie_low_T34Y18;
  wire tie_high_T34Y18;
  wire tie_low_T35Y18;
  wire tie_high_T35Y18;
  wire tie_low_T0Y19;
  wire tie_high_T0Y19;
  wire tie_low_T1Y19;
  wire tie_high_T1Y19;
  wire tie_low_T2Y19;
  wire tie_high_T2Y19;
  wire tie_low_T3Y19;
  wire tie_high_T3Y19;
  wire tie_low_T4Y19;
  wire tie_high_T4Y19;
  wire tie_low_T5Y19;
  wire tie_high_T5Y19;
  wire tie_low_T6Y19;
  wire tie_high_T6Y19;
  wire tie_low_T7Y19;
  wire tie_high_T7Y19;
  wire tie_low_T8Y19;
  wire tie_high_T8Y19;
  wire tie_low_T9Y19;
  wire tie_high_T9Y19;
  wire tie_low_T10Y19;
  wire tie_high_T10Y19;
  wire tie_low_T11Y19;
  wire tie_high_T11Y19;
  wire tie_low_T12Y19;
  wire tie_high_T12Y19;
  wire tie_low_T13Y19;
  wire tie_high_T13Y19;
  wire tie_low_T14Y19;
  wire tie_high_T14Y19;
  wire tie_low_T15Y19;
  wire tie_high_T15Y19;
  wire tie_low_T16Y19;
  wire tie_high_T16Y19;
  wire tie_low_T17Y19;
  wire tie_high_T17Y19;
  wire tie_low_T18Y19;
  wire tie_high_T18Y19;
  wire tie_low_T19Y19;
  wire tie_high_T19Y19;
  wire tie_low_T20Y19;
  wire tie_high_T20Y19;
  wire tie_low_T21Y19;
  wire tie_high_T21Y19;
  wire tie_low_T22Y19;
  wire tie_high_T22Y19;
  wire tie_low_T23Y19;
  wire tie_high_T23Y19;
  wire tie_low_T24Y19;
  wire tie_high_T24Y19;
  wire tie_low_T25Y19;
  wire tie_high_T25Y19;
  wire tie_low_T26Y19;
  wire tie_high_T26Y19;
  wire tie_low_T27Y19;
  wire tie_high_T27Y19;
  wire tie_low_T28Y19;
  wire tie_high_T28Y19;
  wire tie_low_T29Y19;
  wire tie_high_T29Y19;
  wire tie_low_T30Y19;
  wire tie_high_T30Y19;
  wire tie_low_T31Y19;
  wire tie_high_T31Y19;
  wire tie_low_T32Y19;
  wire tie_high_T32Y19;
  wire tie_low_T33Y19;
  wire tie_high_T33Y19;
  wire tie_low_T34Y19;
  wire tie_high_T34Y19;
  wire tie_low_T35Y19;
  wire tie_high_T35Y19;
  wire tie_low_T0Y20;
  wire tie_high_T0Y20;
  wire tie_low_T1Y20;
  wire tie_high_T1Y20;
  wire tie_low_T2Y20;
  wire tie_high_T2Y20;
  wire tie_low_T3Y20;
  wire tie_high_T3Y20;
  wire tie_low_T4Y20;
  wire tie_high_T4Y20;
  wire tie_low_T5Y20;
  wire tie_high_T5Y20;
  wire tie_low_T6Y20;
  wire tie_high_T6Y20;
  wire tie_low_T7Y20;
  wire tie_high_T7Y20;
  wire tie_low_T8Y20;
  wire tie_high_T8Y20;
  wire tie_low_T9Y20;
  wire tie_high_T9Y20;
  wire tie_low_T10Y20;
  wire tie_high_T10Y20;
  wire tie_low_T11Y20;
  wire tie_high_T11Y20;
  wire tie_low_T12Y20;
  wire tie_high_T12Y20;
  wire tie_low_T13Y20;
  wire tie_high_T13Y20;
  wire tie_low_T14Y20;
  wire tie_high_T14Y20;
  wire tie_low_T15Y20;
  wire tie_high_T15Y20;
  wire tie_low_T16Y20;
  wire tie_high_T16Y20;
  wire tie_low_T17Y20;
  wire tie_high_T17Y20;
  wire tie_low_T18Y20;
  wire tie_high_T18Y20;
  wire tie_low_T19Y20;
  wire tie_high_T19Y20;
  wire tie_low_T20Y20;
  wire tie_high_T20Y20;
  wire tie_low_T21Y20;
  wire tie_high_T21Y20;
  wire tie_low_T22Y20;
  wire tie_high_T22Y20;
  wire tie_low_T23Y20;
  wire tie_high_T23Y20;
  wire tie_low_T24Y20;
  wire tie_high_T24Y20;
  wire tie_low_T25Y20;
  wire tie_high_T25Y20;
  wire tie_low_T26Y20;
  wire tie_high_T26Y20;
  wire tie_low_T27Y20;
  wire tie_high_T27Y20;
  wire tie_low_T28Y20;
  wire tie_high_T28Y20;
  wire tie_low_T29Y20;
  wire tie_high_T29Y20;
  wire tie_low_T30Y20;
  wire tie_high_T30Y20;
  wire tie_low_T31Y20;
  wire tie_high_T31Y20;
  wire tie_low_T32Y20;
  wire tie_high_T32Y20;
  wire tie_low_T33Y20;
  wire tie_high_T33Y20;
  wire tie_low_T34Y20;
  wire tie_high_T34Y20;
  wire tie_low_T35Y20;
  wire tie_high_T35Y20;
  wire tie_low_T0Y21;
  wire tie_high_T0Y21;
  wire tie_low_T1Y21;
  wire tie_high_T1Y21;
  wire tie_low_T2Y21;
  wire tie_high_T2Y21;
  wire tie_low_T3Y21;
  wire tie_high_T3Y21;
  wire tie_low_T4Y21;
  wire tie_high_T4Y21;
  wire tie_low_T5Y21;
  wire tie_high_T5Y21;
  wire tie_low_T6Y21;
  wire tie_high_T6Y21;
  wire tie_low_T7Y21;
  wire tie_high_T7Y21;
  wire tie_low_T8Y21;
  wire tie_high_T8Y21;
  wire tie_low_T9Y21;
  wire tie_high_T9Y21;
  wire tie_low_T10Y21;
  wire tie_high_T10Y21;
  wire tie_low_T11Y21;
  wire tie_high_T11Y21;
  wire tie_low_T12Y21;
  wire tie_high_T12Y21;
  wire tie_low_T13Y21;
  wire tie_high_T13Y21;
  wire tie_low_T14Y21;
  wire tie_high_T14Y21;
  wire tie_low_T15Y21;
  wire tie_high_T15Y21;
  wire tie_low_T16Y21;
  wire tie_high_T16Y21;
  wire tie_low_T17Y21;
  wire tie_high_T17Y21;
  wire tie_low_T18Y21;
  wire tie_high_T18Y21;
  wire tie_low_T19Y21;
  wire tie_high_T19Y21;
  wire tie_low_T20Y21;
  wire tie_high_T20Y21;
  wire tie_low_T21Y21;
  wire tie_high_T21Y21;
  wire tie_low_T22Y21;
  wire tie_high_T22Y21;
  wire tie_low_T23Y21;
  wire tie_high_T23Y21;
  wire tie_low_T24Y21;
  wire tie_high_T24Y21;
  wire tie_low_T25Y21;
  wire tie_high_T25Y21;
  wire tie_low_T26Y21;
  wire tie_high_T26Y21;
  wire tie_low_T27Y21;
  wire tie_high_T27Y21;
  wire tie_low_T28Y21;
  wire tie_high_T28Y21;
  wire tie_low_T29Y21;
  wire tie_high_T29Y21;
  wire tie_low_T30Y21;
  wire tie_high_T30Y21;
  wire tie_low_T31Y21;
  wire tie_high_T31Y21;
  wire tie_low_T32Y21;
  wire tie_high_T32Y21;
  wire tie_low_T33Y21;
  wire tie_high_T33Y21;
  wire tie_low_T34Y21;
  wire tie_high_T34Y21;
  wire tie_low_T35Y21;
  wire tie_high_T35Y21;
  wire tie_low_T0Y22;
  wire tie_high_T0Y22;
  wire tie_low_T1Y22;
  wire tie_high_T1Y22;
  wire tie_low_T2Y22;
  wire tie_high_T2Y22;
  wire tie_low_T3Y22;
  wire tie_high_T3Y22;
  wire tie_low_T4Y22;
  wire tie_high_T4Y22;
  wire tie_low_T5Y22;
  wire tie_high_T5Y22;
  wire tie_low_T6Y22;
  wire tie_high_T6Y22;
  wire tie_low_T7Y22;
  wire tie_high_T7Y22;
  wire tie_low_T8Y22;
  wire tie_high_T8Y22;
  wire tie_low_T9Y22;
  wire tie_high_T9Y22;
  wire tie_low_T10Y22;
  wire tie_high_T10Y22;
  wire tie_low_T11Y22;
  wire tie_high_T11Y22;
  wire tie_low_T12Y22;
  wire tie_high_T12Y22;
  wire tie_low_T13Y22;
  wire tie_high_T13Y22;
  wire tie_low_T14Y22;
  wire tie_high_T14Y22;
  wire tie_low_T15Y22;
  wire tie_high_T15Y22;
  wire tie_low_T16Y22;
  wire tie_high_T16Y22;
  wire tie_low_T17Y22;
  wire tie_high_T17Y22;
  wire tie_low_T18Y22;
  wire tie_high_T18Y22;
  wire tie_low_T19Y22;
  wire tie_high_T19Y22;
  wire tie_low_T20Y22;
  wire tie_high_T20Y22;
  wire tie_low_T21Y22;
  wire tie_high_T21Y22;
  wire tie_low_T22Y22;
  wire tie_high_T22Y22;
  wire tie_low_T23Y22;
  wire tie_high_T23Y22;
  wire tie_low_T24Y22;
  wire tie_high_T24Y22;
  wire tie_low_T25Y22;
  wire tie_high_T25Y22;
  wire tie_low_T26Y22;
  wire tie_high_T26Y22;
  wire tie_low_T27Y22;
  wire tie_high_T27Y22;
  wire tie_low_T28Y22;
  wire tie_high_T28Y22;
  wire tie_low_T29Y22;
  wire tie_high_T29Y22;
  wire tie_low_T30Y22;
  wire tie_high_T30Y22;
  wire tie_low_T31Y22;
  wire tie_high_T31Y22;
  wire tie_low_T32Y22;
  wire tie_high_T32Y22;
  wire tie_low_T33Y22;
  wire tie_high_T33Y22;
  wire tie_low_T34Y22;
  wire tie_high_T34Y22;
  wire tie_low_T35Y22;
  wire tie_high_T35Y22;
  wire tie_low_T0Y23;
  wire tie_high_T0Y23;
  wire tie_low_T1Y23;
  wire tie_high_T1Y23;
  wire tie_low_T2Y23;
  wire tie_high_T2Y23;
  wire tie_low_T3Y23;
  wire tie_high_T3Y23;
  wire tie_low_T4Y23;
  wire tie_high_T4Y23;
  wire tie_low_T5Y23;
  wire tie_high_T5Y23;
  wire tie_low_T6Y23;
  wire tie_high_T6Y23;
  wire tie_low_T7Y23;
  wire tie_high_T7Y23;
  wire tie_low_T8Y23;
  wire tie_high_T8Y23;
  wire tie_low_T9Y23;
  wire tie_high_T9Y23;
  wire tie_low_T10Y23;
  wire tie_high_T10Y23;
  wire tie_low_T11Y23;
  wire tie_high_T11Y23;
  wire tie_low_T12Y23;
  wire tie_high_T12Y23;
  wire tie_low_T13Y23;
  wire tie_high_T13Y23;
  wire tie_low_T14Y23;
  wire tie_high_T14Y23;
  wire tie_low_T15Y23;
  wire tie_high_T15Y23;
  wire tie_low_T16Y23;
  wire tie_high_T16Y23;
  wire tie_low_T17Y23;
  wire tie_high_T17Y23;
  wire tie_low_T18Y23;
  wire tie_high_T18Y23;
  wire tie_low_T19Y23;
  wire tie_high_T19Y23;
  wire tie_low_T20Y23;
  wire tie_high_T20Y23;
  wire tie_low_T21Y23;
  wire tie_high_T21Y23;
  wire tie_low_T22Y23;
  wire tie_high_T22Y23;
  wire tie_low_T23Y23;
  wire tie_high_T23Y23;
  wire tie_low_T24Y23;
  wire tie_high_T24Y23;
  wire tie_low_T25Y23;
  wire tie_high_T25Y23;
  wire tie_low_T26Y23;
  wire tie_high_T26Y23;
  wire tie_low_T27Y23;
  wire tie_high_T27Y23;
  wire tie_low_T28Y23;
  wire tie_high_T28Y23;
  wire tie_low_T29Y23;
  wire tie_high_T29Y23;
  wire tie_low_T30Y23;
  wire tie_high_T30Y23;
  wire tie_low_T31Y23;
  wire tie_high_T31Y23;
  wire tie_low_T32Y23;
  wire tie_high_T32Y23;
  wire tie_low_T33Y23;
  wire tie_high_T33Y23;
  wire tie_low_T34Y23;
  wire tie_high_T34Y23;
  wire tie_low_T35Y23;
  wire tie_high_T35Y23;
  wire tie_low_T0Y24;
  wire tie_high_T0Y24;
  wire tie_low_T1Y24;
  wire tie_high_T1Y24;
  wire tie_low_T2Y24;
  wire tie_high_T2Y24;
  wire tie_low_T3Y24;
  wire tie_high_T3Y24;
  wire tie_low_T4Y24;
  wire tie_high_T4Y24;
  wire tie_low_T5Y24;
  wire tie_high_T5Y24;
  wire tie_low_T6Y24;
  wire tie_high_T6Y24;
  wire tie_low_T7Y24;
  wire tie_high_T7Y24;
  wire tie_low_T8Y24;
  wire tie_high_T8Y24;
  wire tie_low_T9Y24;
  wire tie_high_T9Y24;
  wire tie_low_T10Y24;
  wire tie_high_T10Y24;
  wire tie_low_T11Y24;
  wire tie_high_T11Y24;
  wire tie_low_T12Y24;
  wire tie_high_T12Y24;
  wire tie_low_T13Y24;
  wire tie_high_T13Y24;
  wire tie_low_T14Y24;
  wire tie_high_T14Y24;
  wire tie_low_T15Y24;
  wire tie_high_T15Y24;
  wire tie_low_T16Y24;
  wire tie_high_T16Y24;
  wire tie_low_T17Y24;
  wire tie_high_T17Y24;
  wire tie_low_T18Y24;
  wire tie_high_T18Y24;
  wire tie_low_T19Y24;
  wire tie_high_T19Y24;
  wire tie_low_T20Y24;
  wire tie_high_T20Y24;
  wire tie_low_T21Y24;
  wire tie_high_T21Y24;
  wire tie_low_T22Y24;
  wire tie_high_T22Y24;
  wire tie_low_T23Y24;
  wire tie_high_T23Y24;
  wire tie_low_T24Y24;
  wire tie_high_T24Y24;
  wire tie_low_T25Y24;
  wire tie_high_T25Y24;
  wire tie_low_T26Y24;
  wire tie_high_T26Y24;
  wire tie_low_T27Y24;
  wire tie_high_T27Y24;
  wire tie_low_T28Y24;
  wire tie_high_T28Y24;
  wire tie_low_T29Y24;
  wire tie_high_T29Y24;
  wire tie_low_T30Y24;
  wire tie_high_T30Y24;
  wire tie_low_T31Y24;
  wire tie_high_T31Y24;
  wire tie_low_T32Y24;
  wire tie_high_T32Y24;
  wire tie_low_T33Y24;
  wire tie_high_T33Y24;
  wire tie_low_T34Y24;
  wire tie_high_T34Y24;
  wire tie_low_T35Y24;
  wire tie_high_T35Y24;
  wire tie_low_T0Y25;
  wire tie_high_T0Y25;
  wire tie_low_T1Y25;
  wire tie_high_T1Y25;
  wire tie_low_T2Y25;
  wire tie_high_T2Y25;
  wire tie_low_T3Y25;
  wire tie_high_T3Y25;
  wire tie_low_T4Y25;
  wire tie_high_T4Y25;
  wire tie_low_T5Y25;
  wire tie_high_T5Y25;
  wire tie_low_T6Y25;
  wire tie_high_T6Y25;
  wire tie_low_T7Y25;
  wire tie_high_T7Y25;
  wire tie_low_T8Y25;
  wire tie_high_T8Y25;
  wire tie_low_T9Y25;
  wire tie_high_T9Y25;
  wire tie_low_T10Y25;
  wire tie_high_T10Y25;
  wire tie_low_T11Y25;
  wire tie_high_T11Y25;
  wire tie_low_T12Y25;
  wire tie_high_T12Y25;
  wire tie_low_T13Y25;
  wire tie_high_T13Y25;
  wire tie_low_T14Y25;
  wire tie_high_T14Y25;
  wire tie_low_T15Y25;
  wire tie_high_T15Y25;
  wire tie_low_T16Y25;
  wire tie_high_T16Y25;
  wire tie_low_T17Y25;
  wire tie_high_T17Y25;
  wire tie_low_T18Y25;
  wire tie_high_T18Y25;
  wire tie_low_T19Y25;
  wire tie_high_T19Y25;
  wire tie_low_T20Y25;
  wire tie_high_T20Y25;
  wire tie_low_T21Y25;
  wire tie_high_T21Y25;
  wire tie_low_T22Y25;
  wire tie_high_T22Y25;
  wire tie_low_T23Y25;
  wire tie_high_T23Y25;
  wire tie_low_T24Y25;
  wire tie_high_T24Y25;
  wire tie_low_T25Y25;
  wire tie_high_T25Y25;
  wire tie_low_T26Y25;
  wire tie_high_T26Y25;
  wire tie_low_T27Y25;
  wire tie_high_T27Y25;
  wire tie_low_T28Y25;
  wire tie_high_T28Y25;
  wire tie_low_T29Y25;
  wire tie_high_T29Y25;
  wire tie_low_T30Y25;
  wire tie_high_T30Y25;
  wire tie_low_T31Y25;
  wire tie_high_T31Y25;
  wire tie_low_T32Y25;
  wire tie_high_T32Y25;
  wire tie_low_T33Y25;
  wire tie_high_T33Y25;
  wire tie_low_T34Y25;
  wire tie_high_T34Y25;
  wire tie_low_T35Y25;
  wire tie_high_T35Y25;
  wire tie_low_T0Y26;
  wire tie_high_T0Y26;
  wire tie_low_T1Y26;
  wire tie_high_T1Y26;
  wire tie_low_T2Y26;
  wire tie_high_T2Y26;
  wire tie_low_T3Y26;
  wire tie_high_T3Y26;
  wire tie_low_T4Y26;
  wire tie_high_T4Y26;
  wire tie_low_T5Y26;
  wire tie_high_T5Y26;
  wire tie_low_T6Y26;
  wire tie_high_T6Y26;
  wire tie_low_T7Y26;
  wire tie_high_T7Y26;
  wire tie_low_T8Y26;
  wire tie_high_T8Y26;
  wire tie_low_T9Y26;
  wire tie_high_T9Y26;
  wire tie_low_T10Y26;
  wire tie_high_T10Y26;
  wire tie_low_T11Y26;
  wire tie_high_T11Y26;
  wire tie_low_T12Y26;
  wire tie_high_T12Y26;
  wire tie_low_T13Y26;
  wire tie_high_T13Y26;
  wire tie_low_T14Y26;
  wire tie_high_T14Y26;
  wire tie_low_T15Y26;
  wire tie_high_T15Y26;
  wire tie_low_T16Y26;
  wire tie_high_T16Y26;
  wire tie_low_T17Y26;
  wire tie_high_T17Y26;
  wire tie_low_T18Y26;
  wire tie_high_T18Y26;
  wire tie_low_T19Y26;
  wire tie_high_T19Y26;
  wire tie_low_T20Y26;
  wire tie_high_T20Y26;
  wire tie_low_T21Y26;
  wire tie_high_T21Y26;
  wire tie_low_T22Y26;
  wire tie_high_T22Y26;
  wire tie_low_T23Y26;
  wire tie_high_T23Y26;
  wire tie_low_T24Y26;
  wire tie_high_T24Y26;
  wire tie_low_T25Y26;
  wire tie_high_T25Y26;
  wire tie_low_T26Y26;
  wire tie_high_T26Y26;
  wire tie_low_T27Y26;
  wire tie_high_T27Y26;
  wire tie_low_T28Y26;
  wire tie_high_T28Y26;
  wire tie_low_T29Y26;
  wire tie_high_T29Y26;
  wire tie_low_T30Y26;
  wire tie_high_T30Y26;
  wire tie_low_T31Y26;
  wire tie_high_T31Y26;
  wire tie_low_T32Y26;
  wire tie_high_T32Y26;
  wire tie_low_T33Y26;
  wire tie_high_T33Y26;
  wire tie_low_T34Y26;
  wire tie_high_T34Y26;
  wire tie_low_T35Y26;
  wire tie_high_T35Y26;
  wire tie_low_T0Y27;
  wire tie_high_T0Y27;
  wire tie_low_T1Y27;
  wire tie_high_T1Y27;
  wire tie_low_T2Y27;
  wire tie_high_T2Y27;
  wire tie_low_T3Y27;
  wire tie_high_T3Y27;
  wire tie_low_T4Y27;
  wire tie_high_T4Y27;
  wire tie_low_T5Y27;
  wire tie_high_T5Y27;
  wire tie_low_T6Y27;
  wire tie_high_T6Y27;
  wire tie_low_T7Y27;
  wire tie_high_T7Y27;
  wire tie_low_T8Y27;
  wire tie_high_T8Y27;
  wire tie_low_T9Y27;
  wire tie_high_T9Y27;
  wire tie_low_T10Y27;
  wire tie_high_T10Y27;
  wire tie_low_T11Y27;
  wire tie_high_T11Y27;
  wire tie_low_T12Y27;
  wire tie_high_T12Y27;
  wire tie_low_T13Y27;
  wire tie_high_T13Y27;
  wire tie_low_T14Y27;
  wire tie_high_T14Y27;
  wire tie_low_T15Y27;
  wire tie_high_T15Y27;
  wire tie_low_T16Y27;
  wire tie_high_T16Y27;
  wire tie_low_T17Y27;
  wire tie_high_T17Y27;
  wire tie_low_T18Y27;
  wire tie_high_T18Y27;
  wire tie_low_T19Y27;
  wire tie_high_T19Y27;
  wire tie_low_T20Y27;
  wire tie_high_T20Y27;
  wire tie_low_T21Y27;
  wire tie_high_T21Y27;
  wire tie_low_T22Y27;
  wire tie_high_T22Y27;
  wire tie_low_T23Y27;
  wire tie_high_T23Y27;
  wire tie_low_T24Y27;
  wire tie_high_T24Y27;
  wire tie_low_T25Y27;
  wire tie_high_T25Y27;
  wire tie_low_T26Y27;
  wire tie_high_T26Y27;
  wire tie_low_T27Y27;
  wire tie_high_T27Y27;
  wire tie_low_T28Y27;
  wire tie_high_T28Y27;
  wire tie_low_T29Y27;
  wire tie_high_T29Y27;
  wire tie_low_T30Y27;
  wire tie_high_T30Y27;
  wire tie_low_T31Y27;
  wire tie_high_T31Y27;
  wire tie_low_T32Y27;
  wire tie_high_T32Y27;
  wire tie_low_T33Y27;
  wire tie_high_T33Y27;
  wire tie_low_T34Y27;
  wire tie_high_T34Y27;
  wire tie_low_T35Y27;
  wire tie_high_T35Y27;
  wire tie_low_T0Y28;
  wire tie_high_T0Y28;
  wire tie_low_T1Y28;
  wire tie_high_T1Y28;
  wire tie_low_T2Y28;
  wire tie_high_T2Y28;
  wire tie_low_T3Y28;
  wire tie_high_T3Y28;
  wire tie_low_T4Y28;
  wire tie_high_T4Y28;
  wire tie_low_T5Y28;
  wire tie_high_T5Y28;
  wire tie_low_T6Y28;
  wire tie_high_T6Y28;
  wire tie_low_T7Y28;
  wire tie_high_T7Y28;
  wire tie_low_T8Y28;
  wire tie_high_T8Y28;
  wire tie_low_T9Y28;
  wire tie_high_T9Y28;
  wire tie_low_T10Y28;
  wire tie_high_T10Y28;
  wire tie_low_T11Y28;
  wire tie_high_T11Y28;
  wire tie_low_T12Y28;
  wire tie_high_T12Y28;
  wire tie_low_T13Y28;
  wire tie_high_T13Y28;
  wire tie_low_T14Y28;
  wire tie_high_T14Y28;
  wire tie_low_T15Y28;
  wire tie_high_T15Y28;
  wire tie_low_T16Y28;
  wire tie_high_T16Y28;
  wire tie_low_T17Y28;
  wire tie_high_T17Y28;
  wire tie_low_T18Y28;
  wire tie_high_T18Y28;
  wire tie_low_T19Y28;
  wire tie_high_T19Y28;
  wire tie_low_T20Y28;
  wire tie_high_T20Y28;
  wire tie_low_T21Y28;
  wire tie_high_T21Y28;
  wire tie_low_T22Y28;
  wire tie_high_T22Y28;
  wire tie_low_T23Y28;
  wire tie_high_T23Y28;
  wire tie_low_T24Y28;
  wire tie_high_T24Y28;
  wire tie_low_T25Y28;
  wire tie_high_T25Y28;
  wire tie_low_T26Y28;
  wire tie_high_T26Y28;
  wire tie_low_T27Y28;
  wire tie_high_T27Y28;
  wire tie_low_T28Y28;
  wire tie_high_T28Y28;
  wire tie_low_T29Y28;
  wire tie_high_T29Y28;
  wire tie_low_T30Y28;
  wire tie_high_T30Y28;
  wire tie_low_T31Y28;
  wire tie_high_T31Y28;
  wire tie_low_T32Y28;
  wire tie_high_T32Y28;
  wire tie_low_T33Y28;
  wire tie_high_T33Y28;
  wire tie_low_T34Y28;
  wire tie_high_T34Y28;
  wire tie_low_T35Y28;
  wire tie_high_T35Y28;
  wire tie_low_T0Y29;
  wire tie_high_T0Y29;
  wire tie_low_T1Y29;
  wire tie_high_T1Y29;
  wire tie_low_T2Y29;
  wire tie_high_T2Y29;
  wire tie_low_T3Y29;
  wire tie_high_T3Y29;
  wire tie_low_T4Y29;
  wire tie_high_T4Y29;
  wire tie_low_T5Y29;
  wire tie_high_T5Y29;
  wire tie_low_T6Y29;
  wire tie_high_T6Y29;
  wire tie_low_T7Y29;
  wire tie_high_T7Y29;
  wire tie_low_T8Y29;
  wire tie_high_T8Y29;
  wire tie_low_T9Y29;
  wire tie_high_T9Y29;
  wire tie_low_T10Y29;
  wire tie_high_T10Y29;
  wire tie_low_T11Y29;
  wire tie_high_T11Y29;
  wire tie_low_T12Y29;
  wire tie_high_T12Y29;
  wire tie_low_T13Y29;
  wire tie_high_T13Y29;
  wire tie_low_T14Y29;
  wire tie_high_T14Y29;
  wire tie_low_T15Y29;
  wire tie_high_T15Y29;
  wire tie_low_T16Y29;
  wire tie_high_T16Y29;
  wire tie_low_T17Y29;
  wire tie_high_T17Y29;
  wire tie_low_T18Y29;
  wire tie_high_T18Y29;
  wire tie_low_T19Y29;
  wire tie_high_T19Y29;
  wire tie_low_T20Y29;
  wire tie_high_T20Y29;
  wire tie_low_T21Y29;
  wire tie_high_T21Y29;
  wire tie_low_T22Y29;
  wire tie_high_T22Y29;
  wire tie_low_T23Y29;
  wire tie_high_T23Y29;
  wire tie_low_T24Y29;
  wire tie_high_T24Y29;
  wire tie_low_T25Y29;
  wire tie_high_T25Y29;
  wire tie_low_T26Y29;
  wire tie_high_T26Y29;
  wire tie_low_T27Y29;
  wire tie_high_T27Y29;
  wire tie_low_T28Y29;
  wire tie_high_T28Y29;
  wire tie_low_T29Y29;
  wire tie_high_T29Y29;
  wire tie_low_T30Y29;
  wire tie_high_T30Y29;
  wire tie_low_T31Y29;
  wire tie_high_T31Y29;
  wire tie_low_T32Y29;
  wire tie_high_T32Y29;
  wire tie_low_T33Y29;
  wire tie_high_T33Y29;
  wire tie_low_T34Y29;
  wire tie_high_T34Y29;
  wire tie_low_T35Y29;
  wire tie_high_T35Y29;
  wire tie_low_T0Y30;
  wire tie_high_T0Y30;
  wire tie_low_T1Y30;
  wire tie_high_T1Y30;
  wire tie_low_T2Y30;
  wire tie_high_T2Y30;
  wire tie_low_T3Y30;
  wire tie_high_T3Y30;
  wire tie_low_T4Y30;
  wire tie_high_T4Y30;
  wire tie_low_T5Y30;
  wire tie_high_T5Y30;
  wire tie_low_T6Y30;
  wire tie_high_T6Y30;
  wire tie_low_T7Y30;
  wire tie_high_T7Y30;
  wire tie_low_T8Y30;
  wire tie_high_T8Y30;
  wire tie_low_T9Y30;
  wire tie_high_T9Y30;
  wire tie_low_T10Y30;
  wire tie_high_T10Y30;
  wire tie_low_T11Y30;
  wire tie_high_T11Y30;
  wire tie_low_T12Y30;
  wire tie_high_T12Y30;
  wire tie_low_T13Y30;
  wire tie_high_T13Y30;
  wire tie_low_T14Y30;
  wire tie_high_T14Y30;
  wire tie_low_T15Y30;
  wire tie_high_T15Y30;
  wire tie_low_T16Y30;
  wire tie_high_T16Y30;
  wire tie_low_T17Y30;
  wire tie_high_T17Y30;
  wire tie_low_T18Y30;
  wire tie_high_T18Y30;
  wire tie_low_T19Y30;
  wire tie_high_T19Y30;
  wire tie_low_T20Y30;
  wire tie_high_T20Y30;
  wire tie_low_T21Y30;
  wire tie_high_T21Y30;
  wire tie_low_T22Y30;
  wire tie_high_T22Y30;
  wire tie_low_T23Y30;
  wire tie_high_T23Y30;
  wire tie_low_T24Y30;
  wire tie_high_T24Y30;
  wire tie_low_T25Y30;
  wire tie_high_T25Y30;
  wire tie_low_T26Y30;
  wire tie_high_T26Y30;
  wire tie_low_T27Y30;
  wire tie_high_T27Y30;
  wire tie_low_T28Y30;
  wire tie_high_T28Y30;
  wire tie_low_T29Y30;
  wire tie_high_T29Y30;
  wire tie_low_T30Y30;
  wire tie_high_T30Y30;
  wire tie_low_T31Y30;
  wire tie_high_T31Y30;
  wire tie_low_T32Y30;
  wire tie_high_T32Y30;
  wire tie_low_T33Y30;
  wire tie_high_T33Y30;
  wire tie_low_T34Y30;
  wire tie_high_T34Y30;
  wire tie_low_T35Y30;
  wire tie_high_T35Y30;
  wire tie_low_T0Y31;
  wire tie_high_T0Y31;
  wire tie_low_T1Y31;
  wire tie_high_T1Y31;
  wire tie_low_T2Y31;
  wire tie_high_T2Y31;
  wire tie_low_T3Y31;
  wire tie_high_T3Y31;
  wire tie_low_T4Y31;
  wire tie_high_T4Y31;
  wire tie_low_T5Y31;
  wire tie_high_T5Y31;
  wire tie_low_T6Y31;
  wire tie_high_T6Y31;
  wire tie_low_T7Y31;
  wire tie_high_T7Y31;
  wire tie_low_T8Y31;
  wire tie_high_T8Y31;
  wire tie_low_T9Y31;
  wire tie_high_T9Y31;
  wire tie_low_T10Y31;
  wire tie_high_T10Y31;
  wire tie_low_T11Y31;
  wire tie_high_T11Y31;
  wire tie_low_T12Y31;
  wire tie_high_T12Y31;
  wire tie_low_T13Y31;
  wire tie_high_T13Y31;
  wire tie_low_T14Y31;
  wire tie_high_T14Y31;
  wire tie_low_T15Y31;
  wire tie_high_T15Y31;
  wire tie_low_T16Y31;
  wire tie_high_T16Y31;
  wire tie_low_T17Y31;
  wire tie_high_T17Y31;
  wire tie_low_T18Y31;
  wire tie_high_T18Y31;
  wire tie_low_T19Y31;
  wire tie_high_T19Y31;
  wire tie_low_T20Y31;
  wire tie_high_T20Y31;
  wire tie_low_T21Y31;
  wire tie_high_T21Y31;
  wire tie_low_T22Y31;
  wire tie_high_T22Y31;
  wire tie_low_T23Y31;
  wire tie_high_T23Y31;
  wire tie_low_T24Y31;
  wire tie_high_T24Y31;
  wire tie_low_T25Y31;
  wire tie_high_T25Y31;
  wire tie_low_T26Y31;
  wire tie_high_T26Y31;
  wire tie_low_T27Y31;
  wire tie_high_T27Y31;
  wire tie_low_T28Y31;
  wire tie_high_T28Y31;
  wire tie_low_T29Y31;
  wire tie_high_T29Y31;
  wire tie_low_T30Y31;
  wire tie_high_T30Y31;
  wire tie_low_T31Y31;
  wire tie_high_T31Y31;
  wire tie_low_T32Y31;
  wire tie_high_T32Y31;
  wire tie_low_T33Y31;
  wire tie_high_T33Y31;
  wire tie_low_T34Y31;
  wire tie_high_T34Y31;
  wire tie_low_T35Y31;
  wire tie_high_T35Y31;
  wire tie_low_T0Y32;
  wire tie_high_T0Y32;
  wire tie_low_T1Y32;
  wire tie_high_T1Y32;
  wire tie_low_T2Y32;
  wire tie_high_T2Y32;
  wire tie_low_T3Y32;
  wire tie_high_T3Y32;
  wire tie_low_T4Y32;
  wire tie_high_T4Y32;
  wire tie_low_T5Y32;
  wire tie_high_T5Y32;
  wire tie_low_T6Y32;
  wire tie_high_T6Y32;
  wire tie_low_T7Y32;
  wire tie_high_T7Y32;
  wire tie_low_T8Y32;
  wire tie_high_T8Y32;
  wire tie_low_T9Y32;
  wire tie_high_T9Y32;
  wire tie_low_T10Y32;
  wire tie_high_T10Y32;
  wire tie_low_T11Y32;
  wire tie_high_T11Y32;
  wire tie_low_T12Y32;
  wire tie_high_T12Y32;
  wire tie_low_T13Y32;
  wire tie_high_T13Y32;
  wire tie_low_T14Y32;
  wire tie_high_T14Y32;
  wire tie_low_T15Y32;
  wire tie_high_T15Y32;
  wire tie_low_T16Y32;
  wire tie_high_T16Y32;
  wire tie_low_T17Y32;
  wire tie_high_T17Y32;
  wire tie_low_T18Y32;
  wire tie_high_T18Y32;
  wire tie_low_T19Y32;
  wire tie_high_T19Y32;
  wire tie_low_T20Y32;
  wire tie_high_T20Y32;
  wire tie_low_T21Y32;
  wire tie_high_T21Y32;
  wire tie_low_T22Y32;
  wire tie_high_T22Y32;
  wire tie_low_T23Y32;
  wire tie_high_T23Y32;
  wire tie_low_T24Y32;
  wire tie_high_T24Y32;
  wire tie_low_T25Y32;
  wire tie_high_T25Y32;
  wire tie_low_T26Y32;
  wire tie_high_T26Y32;
  wire tie_low_T27Y32;
  wire tie_high_T27Y32;
  wire tie_low_T28Y32;
  wire tie_high_T28Y32;
  wire tie_low_T29Y32;
  wire tie_high_T29Y32;
  wire tie_low_T30Y32;
  wire tie_high_T30Y32;
  wire tie_low_T31Y32;
  wire tie_high_T31Y32;
  wire tie_low_T32Y32;
  wire tie_high_T32Y32;
  wire tie_low_T33Y32;
  wire tie_high_T33Y32;
  wire tie_low_T34Y32;
  wire tie_high_T34Y32;
  wire tie_low_T35Y32;
  wire tie_high_T35Y32;
  wire tie_low_T0Y33;
  wire tie_high_T0Y33;
  wire tie_low_T1Y33;
  wire tie_high_T1Y33;
  wire tie_low_T2Y33;
  wire tie_high_T2Y33;
  wire tie_low_T3Y33;
  wire tie_high_T3Y33;
  wire tie_low_T4Y33;
  wire tie_high_T4Y33;
  wire tie_low_T5Y33;
  wire tie_high_T5Y33;
  wire tie_low_T6Y33;
  wire tie_high_T6Y33;
  wire tie_low_T7Y33;
  wire tie_high_T7Y33;
  wire tie_low_T8Y33;
  wire tie_high_T8Y33;
  wire tie_low_T9Y33;
  wire tie_high_T9Y33;
  wire tie_low_T10Y33;
  wire tie_high_T10Y33;
  wire tie_low_T11Y33;
  wire tie_high_T11Y33;
  wire tie_low_T12Y33;
  wire tie_high_T12Y33;
  wire tie_low_T13Y33;
  wire tie_high_T13Y33;
  wire tie_low_T14Y33;
  wire tie_high_T14Y33;
  wire tie_low_T15Y33;
  wire tie_high_T15Y33;
  wire tie_low_T16Y33;
  wire tie_high_T16Y33;
  wire tie_low_T17Y33;
  wire tie_high_T17Y33;
  wire tie_low_T18Y33;
  wire tie_high_T18Y33;
  wire tie_low_T19Y33;
  wire tie_high_T19Y33;
  wire tie_low_T20Y33;
  wire tie_high_T20Y33;
  wire tie_low_T21Y33;
  wire tie_high_T21Y33;
  wire tie_low_T22Y33;
  wire tie_high_T22Y33;
  wire tie_low_T23Y33;
  wire tie_high_T23Y33;
  wire tie_low_T24Y33;
  wire tie_high_T24Y33;
  wire tie_low_T25Y33;
  wire tie_high_T25Y33;
  wire tie_low_T26Y33;
  wire tie_high_T26Y33;
  wire tie_low_T27Y33;
  wire tie_high_T27Y33;
  wire tie_low_T28Y33;
  wire tie_high_T28Y33;
  wire tie_low_T29Y33;
  wire tie_high_T29Y33;
  wire tie_low_T30Y33;
  wire tie_high_T30Y33;
  wire tie_low_T31Y33;
  wire tie_high_T31Y33;
  wire tie_low_T32Y33;
  wire tie_high_T32Y33;
  wire tie_low_T33Y33;
  wire tie_high_T33Y33;
  wire tie_low_T34Y33;
  wire tie_high_T34Y33;
  wire tie_low_T35Y33;
  wire tie_high_T35Y33;
  wire tie_low_T0Y34;
  wire tie_high_T0Y34;
  wire tie_low_T1Y34;
  wire tie_high_T1Y34;
  wire tie_low_T2Y34;
  wire tie_high_T2Y34;
  wire tie_low_T3Y34;
  wire tie_high_T3Y34;
  wire tie_low_T4Y34;
  wire tie_high_T4Y34;
  wire tie_low_T5Y34;
  wire tie_high_T5Y34;
  wire tie_low_T6Y34;
  wire tie_high_T6Y34;
  wire tie_low_T7Y34;
  wire tie_high_T7Y34;
  wire tie_low_T8Y34;
  wire tie_high_T8Y34;
  wire tie_low_T9Y34;
  wire tie_high_T9Y34;
  wire tie_low_T10Y34;
  wire tie_high_T10Y34;
  wire tie_low_T11Y34;
  wire tie_high_T11Y34;
  wire tie_low_T12Y34;
  wire tie_high_T12Y34;
  wire tie_low_T13Y34;
  wire tie_high_T13Y34;
  wire tie_low_T14Y34;
  wire tie_high_T14Y34;
  wire tie_low_T15Y34;
  wire tie_high_T15Y34;
  wire tie_low_T16Y34;
  wire tie_high_T16Y34;
  wire tie_low_T17Y34;
  wire tie_high_T17Y34;
  wire tie_low_T18Y34;
  wire tie_high_T18Y34;
  wire tie_low_T19Y34;
  wire tie_high_T19Y34;
  wire tie_low_T20Y34;
  wire tie_high_T20Y34;
  wire tie_low_T21Y34;
  wire tie_high_T21Y34;
  wire tie_low_T22Y34;
  wire tie_high_T22Y34;
  wire tie_low_T23Y34;
  wire tie_high_T23Y34;
  wire tie_low_T24Y34;
  wire tie_high_T24Y34;
  wire tie_low_T25Y34;
  wire tie_high_T25Y34;
  wire tie_low_T26Y34;
  wire tie_high_T26Y34;
  wire tie_low_T27Y34;
  wire tie_high_T27Y34;
  wire tie_low_T28Y34;
  wire tie_high_T28Y34;
  wire tie_low_T29Y34;
  wire tie_high_T29Y34;
  wire tie_low_T30Y34;
  wire tie_high_T30Y34;
  wire tie_low_T31Y34;
  wire tie_high_T31Y34;
  wire tie_low_T32Y34;
  wire tie_high_T32Y34;
  wire tie_low_T33Y34;
  wire tie_high_T33Y34;
  wire tie_low_T34Y34;
  wire tie_high_T34Y34;
  wire tie_low_T35Y34;
  wire tie_high_T35Y34;
  wire tie_low_T0Y35;
  wire tie_high_T0Y35;
  wire tie_low_T1Y35;
  wire tie_high_T1Y35;
  wire tie_low_T2Y35;
  wire tie_high_T2Y35;
  wire tie_low_T3Y35;
  wire tie_high_T3Y35;
  wire tie_low_T4Y35;
  wire tie_high_T4Y35;
  wire tie_low_T5Y35;
  wire tie_high_T5Y35;
  wire tie_low_T6Y35;
  wire tie_high_T6Y35;
  wire tie_low_T7Y35;
  wire tie_high_T7Y35;
  wire tie_low_T8Y35;
  wire tie_high_T8Y35;
  wire tie_low_T9Y35;
  wire tie_high_T9Y35;
  wire tie_low_T10Y35;
  wire tie_high_T10Y35;
  wire tie_low_T11Y35;
  wire tie_high_T11Y35;
  wire tie_low_T12Y35;
  wire tie_high_T12Y35;
  wire tie_low_T13Y35;
  wire tie_high_T13Y35;
  wire tie_low_T14Y35;
  wire tie_high_T14Y35;
  wire tie_low_T15Y35;
  wire tie_high_T15Y35;
  wire tie_low_T16Y35;
  wire tie_high_T16Y35;
  wire tie_low_T17Y35;
  wire tie_high_T17Y35;
  wire tie_low_T18Y35;
  wire tie_high_T18Y35;
  wire tie_low_T19Y35;
  wire tie_high_T19Y35;
  wire tie_low_T20Y35;
  wire tie_high_T20Y35;
  wire tie_low_T21Y35;
  wire tie_high_T21Y35;
  wire tie_low_T22Y35;
  wire tie_high_T22Y35;
  wire tie_low_T23Y35;
  wire tie_high_T23Y35;
  wire tie_low_T24Y35;
  wire tie_high_T24Y35;
  wire tie_low_T25Y35;
  wire tie_high_T25Y35;
  wire tie_low_T26Y35;
  wire tie_high_T26Y35;
  wire tie_low_T27Y35;
  wire tie_high_T27Y35;
  wire tie_low_T28Y35;
  wire tie_high_T28Y35;
  wire tie_low_T29Y35;
  wire tie_high_T29Y35;
  wire tie_low_T30Y35;
  wire tie_high_T30Y35;
  wire tie_low_T31Y35;
  wire tie_high_T31Y35;
  wire tie_low_T32Y35;
  wire tie_high_T32Y35;
  wire tie_low_T33Y35;
  wire tie_high_T33Y35;
  wire tie_low_T34Y35;
  wire tie_high_T34Y35;
  wire tie_low_T35Y35;
  wire tie_high_T35Y35;
  wire tie_low_T0Y36;
  wire tie_high_T0Y36;
  wire tie_low_T1Y36;
  wire tie_high_T1Y36;
  wire tie_low_T2Y36;
  wire tie_high_T2Y36;
  wire tie_low_T3Y36;
  wire tie_high_T3Y36;
  wire tie_low_T4Y36;
  wire tie_high_T4Y36;
  wire tie_low_T5Y36;
  wire tie_high_T5Y36;
  wire tie_low_T6Y36;
  wire tie_high_T6Y36;
  wire tie_low_T7Y36;
  wire tie_high_T7Y36;
  wire tie_low_T8Y36;
  wire tie_high_T8Y36;
  wire tie_low_T9Y36;
  wire tie_high_T9Y36;
  wire tie_low_T10Y36;
  wire tie_high_T10Y36;
  wire tie_low_T11Y36;
  wire tie_high_T11Y36;
  wire tie_low_T12Y36;
  wire tie_high_T12Y36;
  wire tie_low_T13Y36;
  wire tie_high_T13Y36;
  wire tie_low_T14Y36;
  wire tie_high_T14Y36;
  wire tie_low_T15Y36;
  wire tie_high_T15Y36;
  wire tie_low_T16Y36;
  wire tie_high_T16Y36;
  wire tie_low_T17Y36;
  wire tie_high_T17Y36;
  wire tie_low_T18Y36;
  wire tie_high_T18Y36;
  wire tie_low_T19Y36;
  wire tie_high_T19Y36;
  wire tie_low_T20Y36;
  wire tie_high_T20Y36;
  wire tie_low_T21Y36;
  wire tie_high_T21Y36;
  wire tie_low_T22Y36;
  wire tie_high_T22Y36;
  wire tie_low_T23Y36;
  wire tie_high_T23Y36;
  wire tie_low_T24Y36;
  wire tie_high_T24Y36;
  wire tie_low_T25Y36;
  wire tie_high_T25Y36;
  wire tie_low_T26Y36;
  wire tie_high_T26Y36;
  wire tie_low_T27Y36;
  wire tie_high_T27Y36;
  wire tie_low_T28Y36;
  wire tie_high_T28Y36;
  wire tie_low_T29Y36;
  wire tie_high_T29Y36;
  wire tie_low_T30Y36;
  wire tie_high_T30Y36;
  wire tie_low_T31Y36;
  wire tie_high_T31Y36;
  wire tie_low_T32Y36;
  wire tie_high_T32Y36;
  wire tie_low_T33Y36;
  wire tie_high_T33Y36;
  wire tie_low_T34Y36;
  wire tie_high_T34Y36;
  wire tie_low_T35Y36;
  wire tie_high_T35Y36;
  wire tie_low_T0Y37;
  wire tie_high_T0Y37;
  wire tie_low_T1Y37;
  wire tie_high_T1Y37;
  wire tie_low_T2Y37;
  wire tie_high_T2Y37;
  wire tie_low_T3Y37;
  wire tie_high_T3Y37;
  wire tie_low_T4Y37;
  wire tie_high_T4Y37;
  wire tie_low_T5Y37;
  wire tie_high_T5Y37;
  wire tie_low_T6Y37;
  wire tie_high_T6Y37;
  wire tie_low_T7Y37;
  wire tie_high_T7Y37;
  wire tie_low_T8Y37;
  wire tie_high_T8Y37;
  wire tie_low_T9Y37;
  wire tie_high_T9Y37;
  wire tie_low_T10Y37;
  wire tie_high_T10Y37;
  wire tie_low_T11Y37;
  wire tie_high_T11Y37;
  wire tie_low_T12Y37;
  wire tie_high_T12Y37;
  wire tie_low_T13Y37;
  wire tie_high_T13Y37;
  wire tie_low_T14Y37;
  wire tie_high_T14Y37;
  wire tie_low_T15Y37;
  wire tie_high_T15Y37;
  wire tie_low_T16Y37;
  wire tie_high_T16Y37;
  wire tie_low_T17Y37;
  wire tie_high_T17Y37;
  wire tie_low_T18Y37;
  wire tie_high_T18Y37;
  wire tie_low_T19Y37;
  wire tie_high_T19Y37;
  wire tie_low_T20Y37;
  wire tie_high_T20Y37;
  wire tie_low_T21Y37;
  wire tie_high_T21Y37;
  wire tie_low_T22Y37;
  wire tie_high_T22Y37;
  wire tie_low_T23Y37;
  wire tie_high_T23Y37;
  wire tie_low_T24Y37;
  wire tie_high_T24Y37;
  wire tie_low_T25Y37;
  wire tie_high_T25Y37;
  wire tie_low_T26Y37;
  wire tie_high_T26Y37;
  wire tie_low_T27Y37;
  wire tie_high_T27Y37;
  wire tie_low_T28Y37;
  wire tie_high_T28Y37;
  wire tie_low_T29Y37;
  wire tie_high_T29Y37;
  wire tie_low_T30Y37;
  wire tie_high_T30Y37;
  wire tie_low_T31Y37;
  wire tie_high_T31Y37;
  wire tie_low_T32Y37;
  wire tie_high_T32Y37;
  wire tie_low_T33Y37;
  wire tie_high_T33Y37;
  wire tie_low_T34Y37;
  wire tie_high_T34Y37;
  wire tie_low_T35Y37;
  wire tie_high_T35Y37;
  wire tie_low_T0Y38;
  wire tie_high_T0Y38;
  wire tie_low_T1Y38;
  wire tie_high_T1Y38;
  wire tie_low_T2Y38;
  wire tie_high_T2Y38;
  wire tie_low_T3Y38;
  wire tie_high_T3Y38;
  wire tie_low_T4Y38;
  wire tie_high_T4Y38;
  wire tie_low_T5Y38;
  wire tie_high_T5Y38;
  wire tie_low_T6Y38;
  wire tie_high_T6Y38;
  wire tie_low_T7Y38;
  wire tie_high_T7Y38;
  wire tie_low_T8Y38;
  wire tie_high_T8Y38;
  wire tie_low_T9Y38;
  wire tie_high_T9Y38;
  wire tie_low_T10Y38;
  wire tie_high_T10Y38;
  wire tie_low_T11Y38;
  wire tie_high_T11Y38;
  wire tie_low_T12Y38;
  wire tie_high_T12Y38;
  wire tie_low_T13Y38;
  wire tie_high_T13Y38;
  wire tie_low_T14Y38;
  wire tie_high_T14Y38;
  wire tie_low_T15Y38;
  wire tie_high_T15Y38;
  wire tie_low_T16Y38;
  wire tie_high_T16Y38;
  wire tie_low_T17Y38;
  wire tie_high_T17Y38;
  wire tie_low_T18Y38;
  wire tie_high_T18Y38;
  wire tie_low_T19Y38;
  wire tie_high_T19Y38;
  wire tie_low_T20Y38;
  wire tie_high_T20Y38;
  wire tie_low_T21Y38;
  wire tie_high_T21Y38;
  wire tie_low_T22Y38;
  wire tie_high_T22Y38;
  wire tie_low_T23Y38;
  wire tie_high_T23Y38;
  wire tie_low_T24Y38;
  wire tie_high_T24Y38;
  wire tie_low_T25Y38;
  wire tie_high_T25Y38;
  wire tie_low_T26Y38;
  wire tie_high_T26Y38;
  wire tie_low_T27Y38;
  wire tie_high_T27Y38;
  wire tie_low_T28Y38;
  wire tie_high_T28Y38;
  wire tie_low_T29Y38;
  wire tie_high_T29Y38;
  wire tie_low_T30Y38;
  wire tie_high_T30Y38;
  wire tie_low_T31Y38;
  wire tie_high_T31Y38;
  wire tie_low_T32Y38;
  wire tie_high_T32Y38;
  wire tie_low_T33Y38;
  wire tie_high_T33Y38;
  wire tie_low_T34Y38;
  wire tie_high_T34Y38;
  wire tie_low_T35Y38;
  wire tie_high_T35Y38;
  wire tie_low_T0Y39;
  wire tie_high_T0Y39;
  wire tie_low_T1Y39;
  wire tie_high_T1Y39;
  wire tie_low_T2Y39;
  wire tie_high_T2Y39;
  wire tie_low_T3Y39;
  wire tie_high_T3Y39;
  wire tie_low_T4Y39;
  wire tie_high_T4Y39;
  wire tie_low_T5Y39;
  wire tie_high_T5Y39;
  wire tie_low_T6Y39;
  wire tie_high_T6Y39;
  wire tie_low_T7Y39;
  wire tie_high_T7Y39;
  wire tie_low_T8Y39;
  wire tie_high_T8Y39;
  wire tie_low_T9Y39;
  wire tie_high_T9Y39;
  wire tie_low_T10Y39;
  wire tie_high_T10Y39;
  wire tie_low_T11Y39;
  wire tie_high_T11Y39;
  wire tie_low_T12Y39;
  wire tie_high_T12Y39;
  wire tie_low_T13Y39;
  wire tie_high_T13Y39;
  wire tie_low_T14Y39;
  wire tie_high_T14Y39;
  wire tie_low_T15Y39;
  wire tie_high_T15Y39;
  wire tie_low_T16Y39;
  wire tie_high_T16Y39;
  wire tie_low_T17Y39;
  wire tie_high_T17Y39;
  wire tie_low_T18Y39;
  wire tie_high_T18Y39;
  wire tie_low_T19Y39;
  wire tie_high_T19Y39;
  wire tie_low_T20Y39;
  wire tie_high_T20Y39;
  wire tie_low_T21Y39;
  wire tie_high_T21Y39;
  wire tie_low_T22Y39;
  wire tie_high_T22Y39;
  wire tie_low_T23Y39;
  wire tie_high_T23Y39;
  wire tie_low_T24Y39;
  wire tie_high_T24Y39;
  wire tie_low_T25Y39;
  wire tie_high_T25Y39;
  wire tie_low_T26Y39;
  wire tie_high_T26Y39;
  wire tie_low_T27Y39;
  wire tie_high_T27Y39;
  wire tie_low_T28Y39;
  wire tie_high_T28Y39;
  wire tie_low_T29Y39;
  wire tie_high_T29Y39;
  wire tie_low_T30Y39;
  wire tie_high_T30Y39;
  wire tie_low_T31Y39;
  wire tie_high_T31Y39;
  wire tie_low_T32Y39;
  wire tie_high_T32Y39;
  wire tie_low_T33Y39;
  wire tie_high_T33Y39;
  wire tie_low_T34Y39;
  wire tie_high_T34Y39;
  wire tie_low_T35Y39;
  wire tie_high_T35Y39;
  wire tie_low_T0Y40;
  wire tie_high_T0Y40;
  wire tie_low_T1Y40;
  wire tie_high_T1Y40;
  wire tie_low_T2Y40;
  wire tie_high_T2Y40;
  wire tie_low_T3Y40;
  wire tie_high_T3Y40;
  wire tie_low_T4Y40;
  wire tie_high_T4Y40;
  wire tie_low_T5Y40;
  wire tie_high_T5Y40;
  wire tie_low_T6Y40;
  wire tie_high_T6Y40;
  wire tie_low_T7Y40;
  wire tie_high_T7Y40;
  wire tie_low_T8Y40;
  wire tie_high_T8Y40;
  wire tie_low_T9Y40;
  wire tie_high_T9Y40;
  wire tie_low_T10Y40;
  wire tie_high_T10Y40;
  wire tie_low_T11Y40;
  wire tie_high_T11Y40;
  wire tie_low_T12Y40;
  wire tie_high_T12Y40;
  wire tie_low_T13Y40;
  wire tie_high_T13Y40;
  wire tie_low_T14Y40;
  wire tie_high_T14Y40;
  wire tie_low_T15Y40;
  wire tie_high_T15Y40;
  wire tie_low_T16Y40;
  wire tie_high_T16Y40;
  wire tie_low_T17Y40;
  wire tie_high_T17Y40;
  wire tie_low_T18Y40;
  wire tie_high_T18Y40;
  wire tie_low_T19Y40;
  wire tie_high_T19Y40;
  wire tie_low_T20Y40;
  wire tie_high_T20Y40;
  wire tie_low_T21Y40;
  wire tie_high_T21Y40;
  wire tie_low_T22Y40;
  wire tie_high_T22Y40;
  wire tie_low_T23Y40;
  wire tie_high_T23Y40;
  wire tie_low_T24Y40;
  wire tie_high_T24Y40;
  wire tie_low_T25Y40;
  wire tie_high_T25Y40;
  wire tie_low_T26Y40;
  wire tie_high_T26Y40;
  wire tie_low_T27Y40;
  wire tie_high_T27Y40;
  wire tie_low_T28Y40;
  wire tie_high_T28Y40;
  wire tie_low_T29Y40;
  wire tie_high_T29Y40;
  wire tie_low_T30Y40;
  wire tie_high_T30Y40;
  wire tie_low_T31Y40;
  wire tie_high_T31Y40;
  wire tie_low_T32Y40;
  wire tie_high_T32Y40;
  wire tie_low_T33Y40;
  wire tie_high_T33Y40;
  wire tie_low_T34Y40;
  wire tie_high_T34Y40;
  wire tie_low_T35Y40;
  wire tie_high_T35Y40;
  wire tie_low_T0Y41;
  wire tie_high_T0Y41;
  wire tie_low_T1Y41;
  wire tie_high_T1Y41;
  wire tie_low_T2Y41;
  wire tie_high_T2Y41;
  wire tie_low_T3Y41;
  wire tie_high_T3Y41;
  wire tie_low_T4Y41;
  wire tie_high_T4Y41;
  wire tie_low_T5Y41;
  wire tie_high_T5Y41;
  wire tie_low_T6Y41;
  wire tie_high_T6Y41;
  wire tie_low_T7Y41;
  wire tie_high_T7Y41;
  wire tie_low_T8Y41;
  wire tie_high_T8Y41;
  wire tie_low_T9Y41;
  wire tie_high_T9Y41;
  wire tie_low_T10Y41;
  wire tie_high_T10Y41;
  wire tie_low_T11Y41;
  wire tie_high_T11Y41;
  wire tie_low_T12Y41;
  wire tie_high_T12Y41;
  wire tie_low_T13Y41;
  wire tie_high_T13Y41;
  wire tie_low_T14Y41;
  wire tie_high_T14Y41;
  wire tie_low_T15Y41;
  wire tie_high_T15Y41;
  wire tie_low_T16Y41;
  wire tie_high_T16Y41;
  wire tie_low_T17Y41;
  wire tie_high_T17Y41;
  wire tie_low_T18Y41;
  wire tie_high_T18Y41;
  wire tie_low_T19Y41;
  wire tie_high_T19Y41;
  wire tie_low_T20Y41;
  wire tie_high_T20Y41;
  wire tie_low_T21Y41;
  wire tie_high_T21Y41;
  wire tie_low_T22Y41;
  wire tie_high_T22Y41;
  wire tie_low_T23Y41;
  wire tie_high_T23Y41;
  wire tie_low_T24Y41;
  wire tie_high_T24Y41;
  wire tie_low_T25Y41;
  wire tie_high_T25Y41;
  wire tie_low_T26Y41;
  wire tie_high_T26Y41;
  wire tie_low_T27Y41;
  wire tie_high_T27Y41;
  wire tie_low_T28Y41;
  wire tie_high_T28Y41;
  wire tie_low_T29Y41;
  wire tie_high_T29Y41;
  wire tie_low_T30Y41;
  wire tie_high_T30Y41;
  wire tie_low_T31Y41;
  wire tie_high_T31Y41;
  wire tie_low_T32Y41;
  wire tie_high_T32Y41;
  wire tie_low_T33Y41;
  wire tie_high_T33Y41;
  wire tie_low_T34Y41;
  wire tie_high_T34Y41;
  wire tie_low_T35Y41;
  wire tie_high_T35Y41;
  wire tie_low_T0Y42;
  wire tie_high_T0Y42;
  wire tie_low_T1Y42;
  wire tie_high_T1Y42;
  wire tie_low_T2Y42;
  wire tie_high_T2Y42;
  wire tie_low_T3Y42;
  wire tie_high_T3Y42;
  wire tie_low_T4Y42;
  wire tie_high_T4Y42;
  wire tie_low_T5Y42;
  wire tie_high_T5Y42;
  wire tie_low_T6Y42;
  wire tie_high_T6Y42;
  wire tie_low_T7Y42;
  wire tie_high_T7Y42;
  wire tie_low_T8Y42;
  wire tie_high_T8Y42;
  wire tie_low_T9Y42;
  wire tie_high_T9Y42;
  wire tie_low_T10Y42;
  wire tie_high_T10Y42;
  wire tie_low_T11Y42;
  wire tie_high_T11Y42;
  wire tie_low_T12Y42;
  wire tie_high_T12Y42;
  wire tie_low_T13Y42;
  wire tie_high_T13Y42;
  wire tie_low_T14Y42;
  wire tie_high_T14Y42;
  wire tie_low_T15Y42;
  wire tie_high_T15Y42;
  wire tie_low_T16Y42;
  wire tie_high_T16Y42;
  wire tie_low_T17Y42;
  wire tie_high_T17Y42;
  wire tie_low_T18Y42;
  wire tie_high_T18Y42;
  wire tie_low_T19Y42;
  wire tie_high_T19Y42;
  wire tie_low_T20Y42;
  wire tie_high_T20Y42;
  wire tie_low_T21Y42;
  wire tie_high_T21Y42;
  wire tie_low_T22Y42;
  wire tie_high_T22Y42;
  wire tie_low_T23Y42;
  wire tie_high_T23Y42;
  wire tie_low_T24Y42;
  wire tie_high_T24Y42;
  wire tie_low_T25Y42;
  wire tie_high_T25Y42;
  wire tie_low_T26Y42;
  wire tie_high_T26Y42;
  wire tie_low_T27Y42;
  wire tie_high_T27Y42;
  wire tie_low_T28Y42;
  wire tie_high_T28Y42;
  wire tie_low_T29Y42;
  wire tie_high_T29Y42;
  wire tie_low_T30Y42;
  wire tie_high_T30Y42;
  wire tie_low_T31Y42;
  wire tie_high_T31Y42;
  wire tie_low_T32Y42;
  wire tie_high_T32Y42;
  wire tie_low_T33Y42;
  wire tie_high_T33Y42;
  wire tie_low_T34Y42;
  wire tie_high_T34Y42;
  wire tie_low_T35Y42;
  wire tie_high_T35Y42;
  wire tie_low_T0Y43;
  wire tie_high_T0Y43;
  wire tie_low_T1Y43;
  wire tie_high_T1Y43;
  wire tie_low_T2Y43;
  wire tie_high_T2Y43;
  wire tie_low_T3Y43;
  wire tie_high_T3Y43;
  wire tie_low_T4Y43;
  wire tie_high_T4Y43;
  wire tie_low_T5Y43;
  wire tie_high_T5Y43;
  wire tie_low_T6Y43;
  wire tie_high_T6Y43;
  wire tie_low_T7Y43;
  wire tie_high_T7Y43;
  wire tie_low_T8Y43;
  wire tie_high_T8Y43;
  wire tie_low_T9Y43;
  wire tie_high_T9Y43;
  wire tie_low_T10Y43;
  wire tie_high_T10Y43;
  wire tie_low_T11Y43;
  wire tie_high_T11Y43;
  wire tie_low_T12Y43;
  wire tie_high_T12Y43;
  wire tie_low_T13Y43;
  wire tie_high_T13Y43;
  wire tie_low_T14Y43;
  wire tie_high_T14Y43;
  wire tie_low_T15Y43;
  wire tie_high_T15Y43;
  wire tie_low_T16Y43;
  wire tie_high_T16Y43;
  wire tie_low_T17Y43;
  wire tie_high_T17Y43;
  wire tie_low_T18Y43;
  wire tie_high_T18Y43;
  wire tie_low_T19Y43;
  wire tie_high_T19Y43;
  wire tie_low_T20Y43;
  wire tie_high_T20Y43;
  wire tie_low_T21Y43;
  wire tie_high_T21Y43;
  wire tie_low_T22Y43;
  wire tie_high_T22Y43;
  wire tie_low_T23Y43;
  wire tie_high_T23Y43;
  wire tie_low_T24Y43;
  wire tie_high_T24Y43;
  wire tie_low_T25Y43;
  wire tie_high_T25Y43;
  wire tie_low_T26Y43;
  wire tie_high_T26Y43;
  wire tie_low_T27Y43;
  wire tie_high_T27Y43;
  wire tie_low_T28Y43;
  wire tie_high_T28Y43;
  wire tie_low_T29Y43;
  wire tie_high_T29Y43;
  wire tie_low_T30Y43;
  wire tie_high_T30Y43;
  wire tie_low_T31Y43;
  wire tie_high_T31Y43;
  wire tie_low_T32Y43;
  wire tie_high_T32Y43;
  wire tie_low_T33Y43;
  wire tie_high_T33Y43;
  wire tie_low_T34Y43;
  wire tie_high_T34Y43;
  wire tie_low_T35Y43;
  wire tie_high_T35Y43;
  wire tie_low_T0Y44;
  wire tie_high_T0Y44;
  wire tie_low_T1Y44;
  wire tie_high_T1Y44;
  wire tie_low_T2Y44;
  wire tie_high_T2Y44;
  wire tie_low_T3Y44;
  wire tie_high_T3Y44;
  wire tie_low_T4Y44;
  wire tie_high_T4Y44;
  wire tie_low_T5Y44;
  wire tie_high_T5Y44;
  wire tie_low_T6Y44;
  wire tie_high_T6Y44;
  wire tie_low_T7Y44;
  wire tie_high_T7Y44;
  wire tie_low_T8Y44;
  wire tie_high_T8Y44;
  wire tie_low_T9Y44;
  wire tie_high_T9Y44;
  wire tie_low_T10Y44;
  wire tie_high_T10Y44;
  wire tie_low_T11Y44;
  wire tie_high_T11Y44;
  wire tie_low_T12Y44;
  wire tie_high_T12Y44;
  wire tie_low_T13Y44;
  wire tie_high_T13Y44;
  wire tie_low_T14Y44;
  wire tie_high_T14Y44;
  wire tie_low_T15Y44;
  wire tie_high_T15Y44;
  wire tie_low_T16Y44;
  wire tie_high_T16Y44;
  wire tie_low_T17Y44;
  wire tie_high_T17Y44;
  wire tie_low_T18Y44;
  wire tie_high_T18Y44;
  wire tie_low_T19Y44;
  wire tie_high_T19Y44;
  wire tie_low_T20Y44;
  wire tie_high_T20Y44;
  wire tie_low_T21Y44;
  wire tie_high_T21Y44;
  wire tie_low_T22Y44;
  wire tie_high_T22Y44;
  wire tie_low_T23Y44;
  wire tie_high_T23Y44;
  wire tie_low_T24Y44;
  wire tie_high_T24Y44;
  wire tie_low_T25Y44;
  wire tie_high_T25Y44;
  wire tie_low_T26Y44;
  wire tie_high_T26Y44;
  wire tie_low_T27Y44;
  wire tie_high_T27Y44;
  wire tie_low_T28Y44;
  wire tie_high_T28Y44;
  wire tie_low_T29Y44;
  wire tie_high_T29Y44;
  wire tie_low_T30Y44;
  wire tie_high_T30Y44;
  wire tie_low_T31Y44;
  wire tie_high_T31Y44;
  wire tie_low_T32Y44;
  wire tie_high_T32Y44;
  wire tie_low_T33Y44;
  wire tie_high_T33Y44;
  wire tie_low_T34Y44;
  wire tie_high_T34Y44;
  wire tie_low_T35Y44;
  wire tie_high_T35Y44;
  wire tie_low_T0Y45;
  wire tie_high_T0Y45;
  wire tie_low_T1Y45;
  wire tie_high_T1Y45;
  wire tie_low_T2Y45;
  wire tie_high_T2Y45;
  wire tie_low_T3Y45;
  wire tie_high_T3Y45;
  wire tie_low_T4Y45;
  wire tie_high_T4Y45;
  wire tie_low_T5Y45;
  wire tie_high_T5Y45;
  wire tie_low_T6Y45;
  wire tie_high_T6Y45;
  wire tie_low_T7Y45;
  wire tie_high_T7Y45;
  wire tie_low_T8Y45;
  wire tie_high_T8Y45;
  wire tie_low_T9Y45;
  wire tie_high_T9Y45;
  wire tie_low_T10Y45;
  wire tie_high_T10Y45;
  wire tie_low_T11Y45;
  wire tie_high_T11Y45;
  wire tie_low_T12Y45;
  wire tie_high_T12Y45;
  wire tie_low_T13Y45;
  wire tie_high_T13Y45;
  wire tie_low_T14Y45;
  wire tie_high_T14Y45;
  wire tie_low_T15Y45;
  wire tie_high_T15Y45;
  wire tie_low_T16Y45;
  wire tie_high_T16Y45;
  wire tie_low_T17Y45;
  wire tie_high_T17Y45;
  wire tie_low_T18Y45;
  wire tie_high_T18Y45;
  wire tie_low_T19Y45;
  wire tie_high_T19Y45;
  wire tie_low_T20Y45;
  wire tie_high_T20Y45;
  wire tie_low_T21Y45;
  wire tie_high_T21Y45;
  wire tie_low_T22Y45;
  wire tie_high_T22Y45;
  wire tie_low_T23Y45;
  wire tie_high_T23Y45;
  wire tie_low_T24Y45;
  wire tie_high_T24Y45;
  wire tie_low_T25Y45;
  wire tie_high_T25Y45;
  wire tie_low_T26Y45;
  wire tie_high_T26Y45;
  wire tie_low_T27Y45;
  wire tie_high_T27Y45;
  wire tie_low_T28Y45;
  wire tie_high_T28Y45;
  wire tie_low_T29Y45;
  wire tie_high_T29Y45;
  wire tie_low_T30Y45;
  wire tie_high_T30Y45;
  wire tie_low_T31Y45;
  wire tie_high_T31Y45;
  wire tie_low_T32Y45;
  wire tie_high_T32Y45;
  wire tie_low_T33Y45;
  wire tie_high_T33Y45;
  wire tie_low_T34Y45;
  wire tie_high_T34Y45;
  wire tie_low_T35Y45;
  wire tie_high_T35Y45;
  wire tie_low_T0Y46;
  wire tie_high_T0Y46;
  wire tie_low_T1Y46;
  wire tie_high_T1Y46;
  wire tie_low_T2Y46;
  wire tie_high_T2Y46;
  wire tie_low_T3Y46;
  wire tie_high_T3Y46;
  wire tie_low_T4Y46;
  wire tie_high_T4Y46;
  wire tie_low_T5Y46;
  wire tie_high_T5Y46;
  wire tie_low_T6Y46;
  wire tie_high_T6Y46;
  wire tie_low_T7Y46;
  wire tie_high_T7Y46;
  wire tie_low_T8Y46;
  wire tie_high_T8Y46;
  wire tie_low_T9Y46;
  wire tie_high_T9Y46;
  wire tie_low_T10Y46;
  wire tie_high_T10Y46;
  wire tie_low_T11Y46;
  wire tie_high_T11Y46;
  wire tie_low_T12Y46;
  wire tie_high_T12Y46;
  wire tie_low_T13Y46;
  wire tie_high_T13Y46;
  wire tie_low_T14Y46;
  wire tie_high_T14Y46;
  wire tie_low_T15Y46;
  wire tie_high_T15Y46;
  wire tie_low_T16Y46;
  wire tie_high_T16Y46;
  wire tie_low_T17Y46;
  wire tie_high_T17Y46;
  wire tie_low_T18Y46;
  wire tie_high_T18Y46;
  wire tie_low_T19Y46;
  wire tie_high_T19Y46;
  wire tie_low_T20Y46;
  wire tie_high_T20Y46;
  wire tie_low_T21Y46;
  wire tie_high_T21Y46;
  wire tie_low_T22Y46;
  wire tie_high_T22Y46;
  wire tie_low_T23Y46;
  wire tie_high_T23Y46;
  wire tie_low_T24Y46;
  wire tie_high_T24Y46;
  wire tie_low_T25Y46;
  wire tie_high_T25Y46;
  wire tie_low_T26Y46;
  wire tie_high_T26Y46;
  wire tie_low_T27Y46;
  wire tie_high_T27Y46;
  wire tie_low_T28Y46;
  wire tie_high_T28Y46;
  wire tie_low_T29Y46;
  wire tie_high_T29Y46;
  wire tie_low_T30Y46;
  wire tie_high_T30Y46;
  wire tie_low_T31Y46;
  wire tie_high_T31Y46;
  wire tie_low_T32Y46;
  wire tie_high_T32Y46;
  wire tie_low_T33Y46;
  wire tie_high_T33Y46;
  wire tie_low_T34Y46;
  wire tie_high_T34Y46;
  wire tie_low_T35Y46;
  wire tie_high_T35Y46;
  wire tie_low_T0Y47;
  wire tie_high_T0Y47;
  wire tie_low_T1Y47;
  wire tie_high_T1Y47;
  wire tie_low_T2Y47;
  wire tie_high_T2Y47;
  wire tie_low_T3Y47;
  wire tie_high_T3Y47;
  wire tie_low_T4Y47;
  wire tie_high_T4Y47;
  wire tie_low_T5Y47;
  wire tie_high_T5Y47;
  wire tie_low_T6Y47;
  wire tie_high_T6Y47;
  wire tie_low_T7Y47;
  wire tie_high_T7Y47;
  wire tie_low_T8Y47;
  wire tie_high_T8Y47;
  wire tie_low_T9Y47;
  wire tie_high_T9Y47;
  wire tie_low_T10Y47;
  wire tie_high_T10Y47;
  wire tie_low_T11Y47;
  wire tie_high_T11Y47;
  wire tie_low_T12Y47;
  wire tie_high_T12Y47;
  wire tie_low_T13Y47;
  wire tie_high_T13Y47;
  wire tie_low_T14Y47;
  wire tie_high_T14Y47;
  wire tie_low_T15Y47;
  wire tie_high_T15Y47;
  wire tie_low_T16Y47;
  wire tie_high_T16Y47;
  wire tie_low_T17Y47;
  wire tie_high_T17Y47;
  wire tie_low_T18Y47;
  wire tie_high_T18Y47;
  wire tie_low_T19Y47;
  wire tie_high_T19Y47;
  wire tie_low_T20Y47;
  wire tie_high_T20Y47;
  wire tie_low_T21Y47;
  wire tie_high_T21Y47;
  wire tie_low_T22Y47;
  wire tie_high_T22Y47;
  wire tie_low_T23Y47;
  wire tie_high_T23Y47;
  wire tie_low_T24Y47;
  wire tie_high_T24Y47;
  wire tie_low_T25Y47;
  wire tie_high_T25Y47;
  wire tie_low_T26Y47;
  wire tie_high_T26Y47;
  wire tie_low_T27Y47;
  wire tie_high_T27Y47;
  wire tie_low_T28Y47;
  wire tie_high_T28Y47;
  wire tie_low_T29Y47;
  wire tie_high_T29Y47;
  wire tie_low_T30Y47;
  wire tie_high_T30Y47;
  wire tie_low_T31Y47;
  wire tie_high_T31Y47;
  wire tie_low_T32Y47;
  wire tie_high_T32Y47;
  wire tie_low_T33Y47;
  wire tie_high_T33Y47;
  wire tie_low_T34Y47;
  wire tie_high_T34Y47;
  wire tie_low_T35Y47;
  wire tie_high_T35Y47;
  wire tie_low_T0Y48;
  wire tie_high_T0Y48;
  wire tie_low_T1Y48;
  wire tie_high_T1Y48;
  wire tie_low_T2Y48;
  wire tie_high_T2Y48;
  wire tie_low_T3Y48;
  wire tie_high_T3Y48;
  wire tie_low_T4Y48;
  wire tie_high_T4Y48;
  wire tie_low_T5Y48;
  wire tie_high_T5Y48;
  wire tie_low_T6Y48;
  wire tie_high_T6Y48;
  wire tie_low_T7Y48;
  wire tie_high_T7Y48;
  wire tie_low_T8Y48;
  wire tie_high_T8Y48;
  wire tie_low_T9Y48;
  wire tie_high_T9Y48;
  wire tie_low_T10Y48;
  wire tie_high_T10Y48;
  wire tie_low_T11Y48;
  wire tie_high_T11Y48;
  wire tie_low_T12Y48;
  wire tie_high_T12Y48;
  wire tie_low_T13Y48;
  wire tie_high_T13Y48;
  wire tie_low_T14Y48;
  wire tie_high_T14Y48;
  wire tie_low_T15Y48;
  wire tie_high_T15Y48;
  wire tie_low_T16Y48;
  wire tie_high_T16Y48;
  wire tie_low_T17Y48;
  wire tie_high_T17Y48;
  wire tie_low_T18Y48;
  wire tie_high_T18Y48;
  wire tie_low_T19Y48;
  wire tie_high_T19Y48;
  wire tie_low_T20Y48;
  wire tie_high_T20Y48;
  wire tie_low_T21Y48;
  wire tie_high_T21Y48;
  wire tie_low_T22Y48;
  wire tie_high_T22Y48;
  wire tie_low_T23Y48;
  wire tie_high_T23Y48;
  wire tie_low_T24Y48;
  wire tie_high_T24Y48;
  wire tie_low_T25Y48;
  wire tie_high_T25Y48;
  wire tie_low_T26Y48;
  wire tie_high_T26Y48;
  wire tie_low_T27Y48;
  wire tie_high_T27Y48;
  wire tie_low_T28Y48;
  wire tie_high_T28Y48;
  wire tie_low_T29Y48;
  wire tie_high_T29Y48;
  wire tie_low_T30Y48;
  wire tie_high_T30Y48;
  wire tie_low_T31Y48;
  wire tie_high_T31Y48;
  wire tie_low_T32Y48;
  wire tie_high_T32Y48;
  wire tie_low_T33Y48;
  wire tie_high_T33Y48;
  wire tie_low_T34Y48;
  wire tie_high_T34Y48;
  wire tie_low_T35Y48;
  wire tie_high_T35Y48;
  wire tie_low_T0Y49;
  wire tie_high_T0Y49;
  wire tie_low_T1Y49;
  wire tie_high_T1Y49;
  wire tie_low_T2Y49;
  wire tie_high_T2Y49;
  wire tie_low_T3Y49;
  wire tie_high_T3Y49;
  wire tie_low_T4Y49;
  wire tie_high_T4Y49;
  wire tie_low_T5Y49;
  wire tie_high_T5Y49;
  wire tie_low_T6Y49;
  wire tie_high_T6Y49;
  wire tie_low_T7Y49;
  wire tie_high_T7Y49;
  wire tie_low_T8Y49;
  wire tie_high_T8Y49;
  wire tie_low_T9Y49;
  wire tie_high_T9Y49;
  wire tie_low_T10Y49;
  wire tie_high_T10Y49;
  wire tie_low_T11Y49;
  wire tie_high_T11Y49;
  wire tie_low_T12Y49;
  wire tie_high_T12Y49;
  wire tie_low_T13Y49;
  wire tie_high_T13Y49;
  wire tie_low_T14Y49;
  wire tie_high_T14Y49;
  wire tie_low_T15Y49;
  wire tie_high_T15Y49;
  wire tie_low_T16Y49;
  wire tie_high_T16Y49;
  wire tie_low_T17Y49;
  wire tie_high_T17Y49;
  wire tie_low_T18Y49;
  wire tie_high_T18Y49;
  wire tie_low_T19Y49;
  wire tie_high_T19Y49;
  wire tie_low_T20Y49;
  wire tie_high_T20Y49;
  wire tie_low_T21Y49;
  wire tie_high_T21Y49;
  wire tie_low_T22Y49;
  wire tie_high_T22Y49;
  wire tie_low_T23Y49;
  wire tie_high_T23Y49;
  wire tie_low_T24Y49;
  wire tie_high_T24Y49;
  wire tie_low_T25Y49;
  wire tie_high_T25Y49;
  wire tie_low_T26Y49;
  wire tie_high_T26Y49;
  wire tie_low_T27Y49;
  wire tie_high_T27Y49;
  wire tie_low_T28Y49;
  wire tie_high_T28Y49;
  wire tie_low_T29Y49;
  wire tie_high_T29Y49;
  wire tie_low_T30Y49;
  wire tie_high_T30Y49;
  wire tie_low_T31Y49;
  wire tie_high_T31Y49;
  wire tie_low_T32Y49;
  wire tie_high_T32Y49;
  wire tie_low_T33Y49;
  wire tie_high_T33Y49;
  wire tie_low_T34Y49;
  wire tie_high_T34Y49;
  wire tie_low_T35Y49;
  wire tie_high_T35Y49;
  wire tie_low_T0Y50;
  wire tie_high_T0Y50;
  wire tie_low_T1Y50;
  wire tie_high_T1Y50;
  wire tie_low_T2Y50;
  wire tie_high_T2Y50;
  wire tie_low_T3Y50;
  wire tie_high_T3Y50;
  wire tie_low_T4Y50;
  wire tie_high_T4Y50;
  wire tie_low_T5Y50;
  wire tie_high_T5Y50;
  wire tie_low_T6Y50;
  wire tie_high_T6Y50;
  wire tie_low_T7Y50;
  wire tie_high_T7Y50;
  wire tie_low_T8Y50;
  wire tie_high_T8Y50;
  wire tie_low_T9Y50;
  wire tie_high_T9Y50;
  wire tie_low_T10Y50;
  wire tie_high_T10Y50;
  wire tie_low_T11Y50;
  wire tie_high_T11Y50;
  wire tie_low_T12Y50;
  wire tie_high_T12Y50;
  wire tie_low_T13Y50;
  wire tie_high_T13Y50;
  wire tie_low_T14Y50;
  wire tie_high_T14Y50;
  wire tie_low_T15Y50;
  wire tie_high_T15Y50;
  wire tie_low_T16Y50;
  wire tie_high_T16Y50;
  wire tie_low_T17Y50;
  wire tie_high_T17Y50;
  wire tie_low_T18Y50;
  wire tie_high_T18Y50;
  wire tie_low_T19Y50;
  wire tie_high_T19Y50;
  wire tie_low_T20Y50;
  wire tie_high_T20Y50;
  wire tie_low_T21Y50;
  wire tie_high_T21Y50;
  wire tie_low_T22Y50;
  wire tie_high_T22Y50;
  wire tie_low_T23Y50;
  wire tie_high_T23Y50;
  wire tie_low_T24Y50;
  wire tie_high_T24Y50;
  wire tie_low_T25Y50;
  wire tie_high_T25Y50;
  wire tie_low_T26Y50;
  wire tie_high_T26Y50;
  wire tie_low_T27Y50;
  wire tie_high_T27Y50;
  wire tie_low_T28Y50;
  wire tie_high_T28Y50;
  wire tie_low_T29Y50;
  wire tie_high_T29Y50;
  wire tie_low_T30Y50;
  wire tie_high_T30Y50;
  wire tie_low_T31Y50;
  wire tie_high_T31Y50;
  wire tie_low_T32Y50;
  wire tie_high_T32Y50;
  wire tie_low_T33Y50;
  wire tie_high_T33Y50;
  wire tie_low_T34Y50;
  wire tie_high_T34Y50;
  wire tie_low_T35Y50;
  wire tie_high_T35Y50;
  wire tie_low_T0Y51;
  wire tie_high_T0Y51;
  wire tie_low_T1Y51;
  wire tie_high_T1Y51;
  wire tie_low_T2Y51;
  wire tie_high_T2Y51;
  wire tie_low_T3Y51;
  wire tie_high_T3Y51;
  wire tie_low_T4Y51;
  wire tie_high_T4Y51;
  wire tie_low_T5Y51;
  wire tie_high_T5Y51;
  wire tie_low_T6Y51;
  wire tie_high_T6Y51;
  wire tie_low_T7Y51;
  wire tie_high_T7Y51;
  wire tie_low_T8Y51;
  wire tie_high_T8Y51;
  wire tie_low_T9Y51;
  wire tie_high_T9Y51;
  wire tie_low_T10Y51;
  wire tie_high_T10Y51;
  wire tie_low_T11Y51;
  wire tie_high_T11Y51;
  wire tie_low_T12Y51;
  wire tie_high_T12Y51;
  wire tie_low_T13Y51;
  wire tie_high_T13Y51;
  wire tie_low_T14Y51;
  wire tie_high_T14Y51;
  wire tie_low_T15Y51;
  wire tie_high_T15Y51;
  wire tie_low_T16Y51;
  wire tie_high_T16Y51;
  wire tie_low_T17Y51;
  wire tie_high_T17Y51;
  wire tie_low_T18Y51;
  wire tie_high_T18Y51;
  wire tie_low_T19Y51;
  wire tie_high_T19Y51;
  wire tie_low_T20Y51;
  wire tie_high_T20Y51;
  wire tie_low_T21Y51;
  wire tie_high_T21Y51;
  wire tie_low_T22Y51;
  wire tie_high_T22Y51;
  wire tie_low_T23Y51;
  wire tie_high_T23Y51;
  wire tie_low_T24Y51;
  wire tie_high_T24Y51;
  wire tie_low_T25Y51;
  wire tie_high_T25Y51;
  wire tie_low_T26Y51;
  wire tie_high_T26Y51;
  wire tie_low_T27Y51;
  wire tie_high_T27Y51;
  wire tie_low_T28Y51;
  wire tie_high_T28Y51;
  wire tie_low_T29Y51;
  wire tie_high_T29Y51;
  wire tie_low_T30Y51;
  wire tie_high_T30Y51;
  wire tie_low_T31Y51;
  wire tie_high_T31Y51;
  wire tie_low_T32Y51;
  wire tie_high_T32Y51;
  wire tie_low_T33Y51;
  wire tie_high_T33Y51;
  wire tie_low_T34Y51;
  wire tie_high_T34Y51;
  wire tie_low_T35Y51;
  wire tie_high_T35Y51;
  wire tie_low_T0Y52;
  wire tie_high_T0Y52;
  wire tie_low_T1Y52;
  wire tie_high_T1Y52;
  wire tie_low_T2Y52;
  wire tie_high_T2Y52;
  wire tie_low_T3Y52;
  wire tie_high_T3Y52;
  wire tie_low_T4Y52;
  wire tie_high_T4Y52;
  wire tie_low_T5Y52;
  wire tie_high_T5Y52;
  wire tie_low_T6Y52;
  wire tie_high_T6Y52;
  wire tie_low_T7Y52;
  wire tie_high_T7Y52;
  wire tie_low_T8Y52;
  wire tie_high_T8Y52;
  wire tie_low_T9Y52;
  wire tie_high_T9Y52;
  wire tie_low_T10Y52;
  wire tie_high_T10Y52;
  wire tie_low_T11Y52;
  wire tie_high_T11Y52;
  wire tie_low_T12Y52;
  wire tie_high_T12Y52;
  wire tie_low_T13Y52;
  wire tie_high_T13Y52;
  wire tie_low_T14Y52;
  wire tie_high_T14Y52;
  wire tie_low_T15Y52;
  wire tie_high_T15Y52;
  wire tie_low_T16Y52;
  wire tie_high_T16Y52;
  wire tie_low_T17Y52;
  wire tie_high_T17Y52;
  wire tie_low_T18Y52;
  wire tie_high_T18Y52;
  wire tie_low_T19Y52;
  wire tie_high_T19Y52;
  wire tie_low_T20Y52;
  wire tie_high_T20Y52;
  wire tie_low_T21Y52;
  wire tie_high_T21Y52;
  wire tie_low_T22Y52;
  wire tie_high_T22Y52;
  wire tie_low_T23Y52;
  wire tie_high_T23Y52;
  wire tie_low_T24Y52;
  wire tie_high_T24Y52;
  wire tie_low_T25Y52;
  wire tie_high_T25Y52;
  wire tie_low_T26Y52;
  wire tie_high_T26Y52;
  wire tie_low_T27Y52;
  wire tie_high_T27Y52;
  wire tie_low_T28Y52;
  wire tie_high_T28Y52;
  wire tie_low_T29Y52;
  wire tie_high_T29Y52;
  wire tie_low_T30Y52;
  wire tie_high_T30Y52;
  wire tie_low_T31Y52;
  wire tie_high_T31Y52;
  wire tie_low_T32Y52;
  wire tie_high_T32Y52;
  wire tie_low_T33Y52;
  wire tie_high_T33Y52;
  wire tie_low_T34Y52;
  wire tie_high_T34Y52;
  wire tie_low_T35Y52;
  wire tie_high_T35Y52;
  wire tie_low_T0Y53;
  wire tie_high_T0Y53;
  wire tie_low_T1Y53;
  wire tie_high_T1Y53;
  wire tie_low_T2Y53;
  wire tie_high_T2Y53;
  wire tie_low_T3Y53;
  wire tie_high_T3Y53;
  wire tie_low_T4Y53;
  wire tie_high_T4Y53;
  wire tie_low_T5Y53;
  wire tie_high_T5Y53;
  wire tie_low_T6Y53;
  wire tie_high_T6Y53;
  wire tie_low_T7Y53;
  wire tie_high_T7Y53;
  wire tie_low_T8Y53;
  wire tie_high_T8Y53;
  wire tie_low_T9Y53;
  wire tie_high_T9Y53;
  wire tie_low_T10Y53;
  wire tie_high_T10Y53;
  wire tie_low_T11Y53;
  wire tie_high_T11Y53;
  wire tie_low_T12Y53;
  wire tie_high_T12Y53;
  wire tie_low_T13Y53;
  wire tie_high_T13Y53;
  wire tie_low_T14Y53;
  wire tie_high_T14Y53;
  wire tie_low_T15Y53;
  wire tie_high_T15Y53;
  wire tie_low_T16Y53;
  wire tie_high_T16Y53;
  wire tie_low_T17Y53;
  wire tie_high_T17Y53;
  wire tie_low_T18Y53;
  wire tie_high_T18Y53;
  wire tie_low_T19Y53;
  wire tie_high_T19Y53;
  wire tie_low_T20Y53;
  wire tie_high_T20Y53;
  wire tie_low_T21Y53;
  wire tie_high_T21Y53;
  wire tie_low_T22Y53;
  wire tie_high_T22Y53;
  wire tie_low_T23Y53;
  wire tie_high_T23Y53;
  wire tie_low_T24Y53;
  wire tie_high_T24Y53;
  wire tie_low_T25Y53;
  wire tie_high_T25Y53;
  wire tie_low_T26Y53;
  wire tie_high_T26Y53;
  wire tie_low_T27Y53;
  wire tie_high_T27Y53;
  wire tie_low_T28Y53;
  wire tie_high_T28Y53;
  wire tie_low_T29Y53;
  wire tie_high_T29Y53;
  wire tie_low_T30Y53;
  wire tie_high_T30Y53;
  wire tie_low_T31Y53;
  wire tie_high_T31Y53;
  wire tie_low_T32Y53;
  wire tie_high_T32Y53;
  wire tie_low_T33Y53;
  wire tie_high_T33Y53;
  wire tie_low_T34Y53;
  wire tie_high_T34Y53;
  wire tie_low_T35Y53;
  wire tie_high_T35Y53;
  wire tie_low_T0Y54;
  wire tie_high_T0Y54;
  wire tie_low_T1Y54;
  wire tie_high_T1Y54;
  wire tie_low_T2Y54;
  wire tie_high_T2Y54;
  wire tie_low_T3Y54;
  wire tie_high_T3Y54;
  wire tie_low_T4Y54;
  wire tie_high_T4Y54;
  wire tie_low_T5Y54;
  wire tie_high_T5Y54;
  wire tie_low_T6Y54;
  wire tie_high_T6Y54;
  wire tie_low_T7Y54;
  wire tie_high_T7Y54;
  wire tie_low_T8Y54;
  wire tie_high_T8Y54;
  wire tie_low_T9Y54;
  wire tie_high_T9Y54;
  wire tie_low_T10Y54;
  wire tie_high_T10Y54;
  wire tie_low_T11Y54;
  wire tie_high_T11Y54;
  wire tie_low_T12Y54;
  wire tie_high_T12Y54;
  wire tie_low_T13Y54;
  wire tie_high_T13Y54;
  wire tie_low_T14Y54;
  wire tie_high_T14Y54;
  wire tie_low_T15Y54;
  wire tie_high_T15Y54;
  wire tie_low_T16Y54;
  wire tie_high_T16Y54;
  wire tie_low_T17Y54;
  wire tie_high_T17Y54;
  wire tie_low_T18Y54;
  wire tie_high_T18Y54;
  wire tie_low_T19Y54;
  wire tie_high_T19Y54;
  wire tie_low_T20Y54;
  wire tie_high_T20Y54;
  wire tie_low_T21Y54;
  wire tie_high_T21Y54;
  wire tie_low_T22Y54;
  wire tie_high_T22Y54;
  wire tie_low_T23Y54;
  wire tie_high_T23Y54;
  wire tie_low_T24Y54;
  wire tie_high_T24Y54;
  wire tie_low_T25Y54;
  wire tie_high_T25Y54;
  wire tie_low_T26Y54;
  wire tie_high_T26Y54;
  wire tie_low_T27Y54;
  wire tie_high_T27Y54;
  wire tie_low_T28Y54;
  wire tie_high_T28Y54;
  wire tie_low_T29Y54;
  wire tie_high_T29Y54;
  wire tie_low_T30Y54;
  wire tie_high_T30Y54;
  wire tie_low_T31Y54;
  wire tie_high_T31Y54;
  wire tie_low_T32Y54;
  wire tie_high_T32Y54;
  wire tie_low_T33Y54;
  wire tie_high_T33Y54;
  wire tie_low_T34Y54;
  wire tie_high_T34Y54;
  wire tie_low_T35Y54;
  wire tie_high_T35Y54;
  wire tie_low_T0Y55;
  wire tie_high_T0Y55;
  wire tie_low_T1Y55;
  wire tie_high_T1Y55;
  wire tie_low_T2Y55;
  wire tie_high_T2Y55;
  wire tie_low_T3Y55;
  wire tie_high_T3Y55;
  wire tie_low_T4Y55;
  wire tie_high_T4Y55;
  wire tie_low_T5Y55;
  wire tie_high_T5Y55;
  wire tie_low_T6Y55;
  wire tie_high_T6Y55;
  wire tie_low_T7Y55;
  wire tie_high_T7Y55;
  wire tie_low_T8Y55;
  wire tie_high_T8Y55;
  wire tie_low_T9Y55;
  wire tie_high_T9Y55;
  wire tie_low_T10Y55;
  wire tie_high_T10Y55;
  wire tie_low_T11Y55;
  wire tie_high_T11Y55;
  wire tie_low_T12Y55;
  wire tie_high_T12Y55;
  wire tie_low_T13Y55;
  wire tie_high_T13Y55;
  wire tie_low_T14Y55;
  wire tie_high_T14Y55;
  wire tie_low_T15Y55;
  wire tie_high_T15Y55;
  wire tie_low_T16Y55;
  wire tie_high_T16Y55;
  wire tie_low_T17Y55;
  wire tie_high_T17Y55;
  wire tie_low_T18Y55;
  wire tie_high_T18Y55;
  wire tie_low_T19Y55;
  wire tie_high_T19Y55;
  wire tie_low_T20Y55;
  wire tie_high_T20Y55;
  wire tie_low_T21Y55;
  wire tie_high_T21Y55;
  wire tie_low_T22Y55;
  wire tie_high_T22Y55;
  wire tie_low_T23Y55;
  wire tie_high_T23Y55;
  wire tie_low_T24Y55;
  wire tie_high_T24Y55;
  wire tie_low_T25Y55;
  wire tie_high_T25Y55;
  wire tie_low_T26Y55;
  wire tie_high_T26Y55;
  wire tie_low_T27Y55;
  wire tie_high_T27Y55;
  wire tie_low_T28Y55;
  wire tie_high_T28Y55;
  wire tie_low_T29Y55;
  wire tie_high_T29Y55;
  wire tie_low_T30Y55;
  wire tie_high_T30Y55;
  wire tie_low_T31Y55;
  wire tie_high_T31Y55;
  wire tie_low_T32Y55;
  wire tie_high_T32Y55;
  wire tie_low_T33Y55;
  wire tie_high_T33Y55;
  wire tie_low_T34Y55;
  wire tie_high_T34Y55;
  wire tie_low_T35Y55;
  wire tie_high_T35Y55;
  wire tie_low_T0Y56;
  wire tie_high_T0Y56;
  wire tie_low_T1Y56;
  wire tie_high_T1Y56;
  wire tie_low_T2Y56;
  wire tie_high_T2Y56;
  wire tie_low_T3Y56;
  wire tie_high_T3Y56;
  wire tie_low_T4Y56;
  wire tie_high_T4Y56;
  wire tie_low_T5Y56;
  wire tie_high_T5Y56;
  wire tie_low_T6Y56;
  wire tie_high_T6Y56;
  wire tie_low_T7Y56;
  wire tie_high_T7Y56;
  wire tie_low_T8Y56;
  wire tie_high_T8Y56;
  wire tie_low_T9Y56;
  wire tie_high_T9Y56;
  wire tie_low_T10Y56;
  wire tie_high_T10Y56;
  wire tie_low_T11Y56;
  wire tie_high_T11Y56;
  wire tie_low_T12Y56;
  wire tie_high_T12Y56;
  wire tie_low_T13Y56;
  wire tie_high_T13Y56;
  wire tie_low_T14Y56;
  wire tie_high_T14Y56;
  wire tie_low_T15Y56;
  wire tie_high_T15Y56;
  wire tie_low_T16Y56;
  wire tie_high_T16Y56;
  wire tie_low_T17Y56;
  wire tie_high_T17Y56;
  wire tie_low_T18Y56;
  wire tie_high_T18Y56;
  wire tie_low_T19Y56;
  wire tie_high_T19Y56;
  wire tie_low_T20Y56;
  wire tie_high_T20Y56;
  wire tie_low_T21Y56;
  wire tie_high_T21Y56;
  wire tie_low_T22Y56;
  wire tie_high_T22Y56;
  wire tie_low_T23Y56;
  wire tie_high_T23Y56;
  wire tie_low_T24Y56;
  wire tie_high_T24Y56;
  wire tie_low_T25Y56;
  wire tie_high_T25Y56;
  wire tie_low_T26Y56;
  wire tie_high_T26Y56;
  wire tie_low_T27Y56;
  wire tie_high_T27Y56;
  wire tie_low_T28Y56;
  wire tie_high_T28Y56;
  wire tie_low_T29Y56;
  wire tie_high_T29Y56;
  wire tie_low_T30Y56;
  wire tie_high_T30Y56;
  wire tie_low_T31Y56;
  wire tie_high_T31Y56;
  wire tie_low_T32Y56;
  wire tie_high_T32Y56;
  wire tie_low_T33Y56;
  wire tie_high_T33Y56;
  wire tie_low_T34Y56;
  wire tie_high_T34Y56;
  wire tie_low_T35Y56;
  wire tie_high_T35Y56;
  wire tie_low_T0Y57;
  wire tie_high_T0Y57;
  wire tie_low_T1Y57;
  wire tie_high_T1Y57;
  wire tie_low_T2Y57;
  wire tie_high_T2Y57;
  wire tie_low_T3Y57;
  wire tie_high_T3Y57;
  wire tie_low_T4Y57;
  wire tie_high_T4Y57;
  wire tie_low_T5Y57;
  wire tie_high_T5Y57;
  wire tie_low_T6Y57;
  wire tie_high_T6Y57;
  wire tie_low_T7Y57;
  wire tie_high_T7Y57;
  wire tie_low_T8Y57;
  wire tie_high_T8Y57;
  wire tie_low_T9Y57;
  wire tie_high_T9Y57;
  wire tie_low_T10Y57;
  wire tie_high_T10Y57;
  wire tie_low_T11Y57;
  wire tie_high_T11Y57;
  wire tie_low_T12Y57;
  wire tie_high_T12Y57;
  wire tie_low_T13Y57;
  wire tie_high_T13Y57;
  wire tie_low_T14Y57;
  wire tie_high_T14Y57;
  wire tie_low_T15Y57;
  wire tie_high_T15Y57;
  wire tie_low_T16Y57;
  wire tie_high_T16Y57;
  wire tie_low_T17Y57;
  wire tie_high_T17Y57;
  wire tie_low_T18Y57;
  wire tie_high_T18Y57;
  wire tie_low_T19Y57;
  wire tie_high_T19Y57;
  wire tie_low_T20Y57;
  wire tie_high_T20Y57;
  wire tie_low_T21Y57;
  wire tie_high_T21Y57;
  wire tie_low_T22Y57;
  wire tie_high_T22Y57;
  wire tie_low_T23Y57;
  wire tie_high_T23Y57;
  wire tie_low_T24Y57;
  wire tie_high_T24Y57;
  wire tie_low_T25Y57;
  wire tie_high_T25Y57;
  wire tie_low_T26Y57;
  wire tie_high_T26Y57;
  wire tie_low_T27Y57;
  wire tie_high_T27Y57;
  wire tie_low_T28Y57;
  wire tie_high_T28Y57;
  wire tie_low_T29Y57;
  wire tie_high_T29Y57;
  wire tie_low_T30Y57;
  wire tie_high_T30Y57;
  wire tie_low_T31Y57;
  wire tie_high_T31Y57;
  wire tie_low_T32Y57;
  wire tie_high_T32Y57;
  wire tie_low_T33Y57;
  wire tie_high_T33Y57;
  wire tie_low_T34Y57;
  wire tie_high_T34Y57;
  wire tie_low_T35Y57;
  wire tie_high_T35Y57;
  wire tie_low_T0Y58;
  wire tie_high_T0Y58;
  wire tie_low_T1Y58;
  wire tie_high_T1Y58;
  wire tie_low_T2Y58;
  wire tie_high_T2Y58;
  wire tie_low_T3Y58;
  wire tie_high_T3Y58;
  wire tie_low_T4Y58;
  wire tie_high_T4Y58;
  wire tie_low_T5Y58;
  wire tie_high_T5Y58;
  wire tie_low_T6Y58;
  wire tie_high_T6Y58;
  wire tie_low_T7Y58;
  wire tie_high_T7Y58;
  wire tie_low_T8Y58;
  wire tie_high_T8Y58;
  wire tie_low_T9Y58;
  wire tie_high_T9Y58;
  wire tie_low_T10Y58;
  wire tie_high_T10Y58;
  wire tie_low_T11Y58;
  wire tie_high_T11Y58;
  wire tie_low_T12Y58;
  wire tie_high_T12Y58;
  wire tie_low_T13Y58;
  wire tie_high_T13Y58;
  wire tie_low_T14Y58;
  wire tie_high_T14Y58;
  wire tie_low_T15Y58;
  wire tie_high_T15Y58;
  wire tie_low_T16Y58;
  wire tie_high_T16Y58;
  wire tie_low_T17Y58;
  wire tie_high_T17Y58;
  wire tie_low_T18Y58;
  wire tie_high_T18Y58;
  wire tie_low_T19Y58;
  wire tie_high_T19Y58;
  wire tie_low_T20Y58;
  wire tie_high_T20Y58;
  wire tie_low_T21Y58;
  wire tie_high_T21Y58;
  wire tie_low_T22Y58;
  wire tie_high_T22Y58;
  wire tie_low_T23Y58;
  wire tie_high_T23Y58;
  wire tie_low_T24Y58;
  wire tie_high_T24Y58;
  wire tie_low_T25Y58;
  wire tie_high_T25Y58;
  wire tie_low_T26Y58;
  wire tie_high_T26Y58;
  wire tie_low_T27Y58;
  wire tie_high_T27Y58;
  wire tie_low_T28Y58;
  wire tie_high_T28Y58;
  wire tie_low_T29Y58;
  wire tie_high_T29Y58;
  wire tie_low_T30Y58;
  wire tie_high_T30Y58;
  wire tie_low_T31Y58;
  wire tie_high_T31Y58;
  wire tie_low_T32Y58;
  wire tie_high_T32Y58;
  wire tie_low_T33Y58;
  wire tie_high_T33Y58;
  wire tie_low_T34Y58;
  wire tie_high_T34Y58;
  wire tie_low_T35Y58;
  wire tie_high_T35Y58;
  wire tie_low_T0Y59;
  wire tie_high_T0Y59;
  wire tie_low_T1Y59;
  wire tie_high_T1Y59;
  wire tie_low_T2Y59;
  wire tie_high_T2Y59;
  wire tie_low_T3Y59;
  wire tie_high_T3Y59;
  wire tie_low_T4Y59;
  wire tie_high_T4Y59;
  wire tie_low_T5Y59;
  wire tie_high_T5Y59;
  wire tie_low_T6Y59;
  wire tie_high_T6Y59;
  wire tie_low_T7Y59;
  wire tie_high_T7Y59;
  wire tie_low_T8Y59;
  wire tie_high_T8Y59;
  wire tie_low_T9Y59;
  wire tie_high_T9Y59;
  wire tie_low_T10Y59;
  wire tie_high_T10Y59;
  wire tie_low_T11Y59;
  wire tie_high_T11Y59;
  wire tie_low_T12Y59;
  wire tie_high_T12Y59;
  wire tie_low_T13Y59;
  wire tie_high_T13Y59;
  wire tie_low_T14Y59;
  wire tie_high_T14Y59;
  wire tie_low_T15Y59;
  wire tie_high_T15Y59;
  wire tie_low_T16Y59;
  wire tie_high_T16Y59;
  wire tie_low_T17Y59;
  wire tie_high_T17Y59;
  wire tie_low_T18Y59;
  wire tie_high_T18Y59;
  wire tie_low_T19Y59;
  wire tie_high_T19Y59;
  wire tie_low_T20Y59;
  wire tie_high_T20Y59;
  wire tie_low_T21Y59;
  wire tie_high_T21Y59;
  wire tie_low_T22Y59;
  wire tie_high_T22Y59;
  wire tie_low_T23Y59;
  wire tie_high_T23Y59;
  wire tie_low_T24Y59;
  wire tie_high_T24Y59;
  wire tie_low_T25Y59;
  wire tie_high_T25Y59;
  wire tie_low_T26Y59;
  wire tie_high_T26Y59;
  wire tie_low_T27Y59;
  wire tie_high_T27Y59;
  wire tie_low_T28Y59;
  wire tie_high_T28Y59;
  wire tie_low_T29Y59;
  wire tie_high_T29Y59;
  wire tie_low_T30Y59;
  wire tie_high_T30Y59;
  wire tie_low_T31Y59;
  wire tie_high_T31Y59;
  wire tie_low_T32Y59;
  wire tie_high_T32Y59;
  wire tie_low_T33Y59;
  wire tie_high_T33Y59;
  wire tie_low_T34Y59;
  wire tie_high_T34Y59;
  wire tie_low_T35Y59;
  wire tie_high_T35Y59;
  wire tie_low_T0Y60;
  wire tie_high_T0Y60;
  wire tie_low_T1Y60;
  wire tie_high_T1Y60;
  wire tie_low_T2Y60;
  wire tie_high_T2Y60;
  wire tie_low_T3Y60;
  wire tie_high_T3Y60;
  wire tie_low_T4Y60;
  wire tie_high_T4Y60;
  wire tie_low_T5Y60;
  wire tie_high_T5Y60;
  wire tie_low_T6Y60;
  wire tie_high_T6Y60;
  wire tie_low_T7Y60;
  wire tie_high_T7Y60;
  wire tie_low_T8Y60;
  wire tie_high_T8Y60;
  wire tie_low_T9Y60;
  wire tie_high_T9Y60;
  wire tie_low_T10Y60;
  wire tie_high_T10Y60;
  wire tie_low_T11Y60;
  wire tie_high_T11Y60;
  wire tie_low_T12Y60;
  wire tie_high_T12Y60;
  wire tie_low_T13Y60;
  wire tie_high_T13Y60;
  wire tie_low_T14Y60;
  wire tie_high_T14Y60;
  wire tie_low_T15Y60;
  wire tie_high_T15Y60;
  wire tie_low_T16Y60;
  wire tie_high_T16Y60;
  wire tie_low_T17Y60;
  wire tie_high_T17Y60;
  wire tie_low_T18Y60;
  wire tie_high_T18Y60;
  wire tie_low_T19Y60;
  wire tie_high_T19Y60;
  wire tie_low_T20Y60;
  wire tie_high_T20Y60;
  wire tie_low_T21Y60;
  wire tie_high_T21Y60;
  wire tie_low_T22Y60;
  wire tie_high_T22Y60;
  wire tie_low_T23Y60;
  wire tie_high_T23Y60;
  wire tie_low_T24Y60;
  wire tie_high_T24Y60;
  wire tie_low_T25Y60;
  wire tie_high_T25Y60;
  wire tie_low_T26Y60;
  wire tie_high_T26Y60;
  wire tie_low_T27Y60;
  wire tie_high_T27Y60;
  wire tie_low_T28Y60;
  wire tie_high_T28Y60;
  wire tie_low_T29Y60;
  wire tie_high_T29Y60;
  wire tie_low_T30Y60;
  wire tie_high_T30Y60;
  wire tie_low_T31Y60;
  wire tie_high_T31Y60;
  wire tie_low_T32Y60;
  wire tie_high_T32Y60;
  wire tie_low_T33Y60;
  wire tie_high_T33Y60;
  wire tie_low_T34Y60;
  wire tie_high_T34Y60;
  wire tie_low_T35Y60;
  wire tie_high_T35Y60;
  wire tie_low_T0Y61;
  wire tie_high_T0Y61;
  wire tie_low_T1Y61;
  wire tie_high_T1Y61;
  wire tie_low_T2Y61;
  wire tie_high_T2Y61;
  wire tie_low_T3Y61;
  wire tie_high_T3Y61;
  wire tie_low_T4Y61;
  wire tie_high_T4Y61;
  wire tie_low_T5Y61;
  wire tie_high_T5Y61;
  wire tie_low_T6Y61;
  wire tie_high_T6Y61;
  wire tie_low_T7Y61;
  wire tie_high_T7Y61;
  wire tie_low_T8Y61;
  wire tie_high_T8Y61;
  wire tie_low_T9Y61;
  wire tie_high_T9Y61;
  wire tie_low_T10Y61;
  wire tie_high_T10Y61;
  wire tie_low_T11Y61;
  wire tie_high_T11Y61;
  wire tie_low_T12Y61;
  wire tie_high_T12Y61;
  wire tie_low_T13Y61;
  wire tie_high_T13Y61;
  wire tie_low_T14Y61;
  wire tie_high_T14Y61;
  wire tie_low_T15Y61;
  wire tie_high_T15Y61;
  wire tie_low_T16Y61;
  wire tie_high_T16Y61;
  wire tie_low_T17Y61;
  wire tie_high_T17Y61;
  wire tie_low_T18Y61;
  wire tie_high_T18Y61;
  wire tie_low_T19Y61;
  wire tie_high_T19Y61;
  wire tie_low_T20Y61;
  wire tie_high_T20Y61;
  wire tie_low_T21Y61;
  wire tie_high_T21Y61;
  wire tie_low_T22Y61;
  wire tie_high_T22Y61;
  wire tie_low_T23Y61;
  wire tie_high_T23Y61;
  wire tie_low_T24Y61;
  wire tie_high_T24Y61;
  wire tie_low_T25Y61;
  wire tie_high_T25Y61;
  wire tie_low_T26Y61;
  wire tie_high_T26Y61;
  wire tie_low_T27Y61;
  wire tie_high_T27Y61;
  wire tie_low_T28Y61;
  wire tie_high_T28Y61;
  wire tie_low_T29Y61;
  wire tie_high_T29Y61;
  wire tie_low_T30Y61;
  wire tie_high_T30Y61;
  wire tie_low_T31Y61;
  wire tie_high_T31Y61;
  wire tie_low_T32Y61;
  wire tie_high_T32Y61;
  wire tie_low_T33Y61;
  wire tie_high_T33Y61;
  wire tie_low_T34Y61;
  wire tie_high_T34Y61;
  wire tie_low_T35Y61;
  wire tie_high_T35Y61;
  wire tie_low_T0Y62;
  wire tie_high_T0Y62;
  wire tie_low_T1Y62;
  wire tie_high_T1Y62;
  wire tie_low_T2Y62;
  wire tie_high_T2Y62;
  wire tie_low_T3Y62;
  wire tie_high_T3Y62;
  wire tie_low_T4Y62;
  wire tie_high_T4Y62;
  wire tie_low_T5Y62;
  wire tie_high_T5Y62;
  wire tie_low_T6Y62;
  wire tie_high_T6Y62;
  wire tie_low_T7Y62;
  wire tie_high_T7Y62;
  wire tie_low_T8Y62;
  wire tie_high_T8Y62;
  wire tie_low_T9Y62;
  wire tie_high_T9Y62;
  wire tie_low_T10Y62;
  wire tie_high_T10Y62;
  wire tie_low_T11Y62;
  wire tie_high_T11Y62;
  wire tie_low_T12Y62;
  wire tie_high_T12Y62;
  wire tie_low_T13Y62;
  wire tie_high_T13Y62;
  wire tie_low_T14Y62;
  wire tie_high_T14Y62;
  wire tie_low_T15Y62;
  wire tie_high_T15Y62;
  wire tie_low_T16Y62;
  wire tie_high_T16Y62;
  wire tie_low_T17Y62;
  wire tie_high_T17Y62;
  wire tie_low_T18Y62;
  wire tie_high_T18Y62;
  wire tie_low_T19Y62;
  wire tie_high_T19Y62;
  wire tie_low_T20Y62;
  wire tie_high_T20Y62;
  wire tie_low_T21Y62;
  wire tie_high_T21Y62;
  wire tie_low_T22Y62;
  wire tie_high_T22Y62;
  wire tie_low_T23Y62;
  wire tie_high_T23Y62;
  wire tie_low_T24Y62;
  wire tie_high_T24Y62;
  wire tie_low_T25Y62;
  wire tie_high_T25Y62;
  wire tie_low_T26Y62;
  wire tie_high_T26Y62;
  wire tie_low_T27Y62;
  wire tie_high_T27Y62;
  wire tie_low_T28Y62;
  wire tie_high_T28Y62;
  wire tie_low_T29Y62;
  wire tie_high_T29Y62;
  wire tie_low_T30Y62;
  wire tie_high_T30Y62;
  wire tie_low_T31Y62;
  wire tie_high_T31Y62;
  wire tie_low_T32Y62;
  wire tie_high_T32Y62;
  wire tie_low_T33Y62;
  wire tie_high_T33Y62;
  wire tie_low_T34Y62;
  wire tie_high_T34Y62;
  wire tie_low_T35Y62;
  wire tie_high_T35Y62;
  wire tie_low_T0Y63;
  wire tie_high_T0Y63;
  wire tie_low_T1Y63;
  wire tie_high_T1Y63;
  wire tie_low_T2Y63;
  wire tie_high_T2Y63;
  wire tie_low_T3Y63;
  wire tie_high_T3Y63;
  wire tie_low_T4Y63;
  wire tie_high_T4Y63;
  wire tie_low_T5Y63;
  wire tie_high_T5Y63;
  wire tie_low_T6Y63;
  wire tie_high_T6Y63;
  wire tie_low_T7Y63;
  wire tie_high_T7Y63;
  wire tie_low_T8Y63;
  wire tie_high_T8Y63;
  wire tie_low_T9Y63;
  wire tie_high_T9Y63;
  wire tie_low_T10Y63;
  wire tie_high_T10Y63;
  wire tie_low_T11Y63;
  wire tie_high_T11Y63;
  wire tie_low_T12Y63;
  wire tie_high_T12Y63;
  wire tie_low_T13Y63;
  wire tie_high_T13Y63;
  wire tie_low_T14Y63;
  wire tie_high_T14Y63;
  wire tie_low_T15Y63;
  wire tie_high_T15Y63;
  wire tie_low_T16Y63;
  wire tie_high_T16Y63;
  wire tie_low_T17Y63;
  wire tie_high_T17Y63;
  wire tie_low_T18Y63;
  wire tie_high_T18Y63;
  wire tie_low_T19Y63;
  wire tie_high_T19Y63;
  wire tie_low_T20Y63;
  wire tie_high_T20Y63;
  wire tie_low_T21Y63;
  wire tie_high_T21Y63;
  wire tie_low_T22Y63;
  wire tie_high_T22Y63;
  wire tie_low_T23Y63;
  wire tie_high_T23Y63;
  wire tie_low_T24Y63;
  wire tie_high_T24Y63;
  wire tie_low_T25Y63;
  wire tie_high_T25Y63;
  wire tie_low_T26Y63;
  wire tie_high_T26Y63;
  wire tie_low_T27Y63;
  wire tie_high_T27Y63;
  wire tie_low_T28Y63;
  wire tie_high_T28Y63;
  wire tie_low_T29Y63;
  wire tie_high_T29Y63;
  wire tie_low_T30Y63;
  wire tie_high_T30Y63;
  wire tie_low_T31Y63;
  wire tie_high_T31Y63;
  wire tie_low_T32Y63;
  wire tie_high_T32Y63;
  wire tie_low_T33Y63;
  wire tie_high_T33Y63;
  wire tie_low_T34Y63;
  wire tie_high_T34Y63;
  wire tie_low_T35Y63;
  wire tie_high_T35Y63;
  wire tie_low_T0Y64;
  wire tie_high_T0Y64;
  wire tie_low_T1Y64;
  wire tie_high_T1Y64;
  wire tie_low_T2Y64;
  wire tie_high_T2Y64;
  wire tie_low_T3Y64;
  wire tie_high_T3Y64;
  wire tie_low_T4Y64;
  wire tie_high_T4Y64;
  wire tie_low_T5Y64;
  wire tie_high_T5Y64;
  wire tie_low_T6Y64;
  wire tie_high_T6Y64;
  wire tie_low_T7Y64;
  wire tie_high_T7Y64;
  wire tie_low_T8Y64;
  wire tie_high_T8Y64;
  wire tie_low_T9Y64;
  wire tie_high_T9Y64;
  wire tie_low_T10Y64;
  wire tie_high_T10Y64;
  wire tie_low_T11Y64;
  wire tie_high_T11Y64;
  wire tie_low_T12Y64;
  wire tie_high_T12Y64;
  wire tie_low_T13Y64;
  wire tie_high_T13Y64;
  wire tie_low_T14Y64;
  wire tie_high_T14Y64;
  wire tie_low_T15Y64;
  wire tie_high_T15Y64;
  wire tie_low_T16Y64;
  wire tie_high_T16Y64;
  wire tie_low_T17Y64;
  wire tie_high_T17Y64;
  wire tie_low_T18Y64;
  wire tie_high_T18Y64;
  wire tie_low_T19Y64;
  wire tie_high_T19Y64;
  wire tie_low_T20Y64;
  wire tie_high_T20Y64;
  wire tie_low_T21Y64;
  wire tie_high_T21Y64;
  wire tie_low_T22Y64;
  wire tie_high_T22Y64;
  wire tie_low_T23Y64;
  wire tie_high_T23Y64;
  wire tie_low_T24Y64;
  wire tie_high_T24Y64;
  wire tie_low_T25Y64;
  wire tie_high_T25Y64;
  wire tie_low_T26Y64;
  wire tie_high_T26Y64;
  wire tie_low_T27Y64;
  wire tie_high_T27Y64;
  wire tie_low_T28Y64;
  wire tie_high_T28Y64;
  wire tie_low_T29Y64;
  wire tie_high_T29Y64;
  wire tie_low_T30Y64;
  wire tie_high_T30Y64;
  wire tie_low_T31Y64;
  wire tie_high_T31Y64;
  wire tie_low_T32Y64;
  wire tie_high_T32Y64;
  wire tie_low_T33Y64;
  wire tie_high_T33Y64;
  wire tie_low_T34Y64;
  wire tie_high_T34Y64;
  wire tie_low_T35Y64;
  wire tie_high_T35Y64;
  wire tie_low_T0Y65;
  wire tie_high_T0Y65;
  wire tie_low_T1Y65;
  wire tie_high_T1Y65;
  wire tie_low_T2Y65;
  wire tie_high_T2Y65;
  wire tie_low_T3Y65;
  wire tie_high_T3Y65;
  wire tie_low_T4Y65;
  wire tie_high_T4Y65;
  wire tie_low_T5Y65;
  wire tie_high_T5Y65;
  wire tie_low_T6Y65;
  wire tie_high_T6Y65;
  wire tie_low_T7Y65;
  wire tie_high_T7Y65;
  wire tie_low_T8Y65;
  wire tie_high_T8Y65;
  wire tie_low_T9Y65;
  wire tie_high_T9Y65;
  wire tie_low_T10Y65;
  wire tie_high_T10Y65;
  wire tie_low_T11Y65;
  wire tie_high_T11Y65;
  wire tie_low_T12Y65;
  wire tie_high_T12Y65;
  wire tie_low_T13Y65;
  wire tie_high_T13Y65;
  wire tie_low_T14Y65;
  wire tie_high_T14Y65;
  wire tie_low_T15Y65;
  wire tie_high_T15Y65;
  wire tie_low_T16Y65;
  wire tie_high_T16Y65;
  wire tie_low_T17Y65;
  wire tie_high_T17Y65;
  wire tie_low_T18Y65;
  wire tie_high_T18Y65;
  wire tie_low_T19Y65;
  wire tie_high_T19Y65;
  wire tie_low_T20Y65;
  wire tie_high_T20Y65;
  wire tie_low_T21Y65;
  wire tie_high_T21Y65;
  wire tie_low_T22Y65;
  wire tie_high_T22Y65;
  wire tie_low_T23Y65;
  wire tie_high_T23Y65;
  wire tie_low_T24Y65;
  wire tie_high_T24Y65;
  wire tie_low_T25Y65;
  wire tie_high_T25Y65;
  wire tie_low_T26Y65;
  wire tie_high_T26Y65;
  wire tie_low_T27Y65;
  wire tie_high_T27Y65;
  wire tie_low_T28Y65;
  wire tie_high_T28Y65;
  wire tie_low_T29Y65;
  wire tie_high_T29Y65;
  wire tie_low_T30Y65;
  wire tie_high_T30Y65;
  wire tie_low_T31Y65;
  wire tie_high_T31Y65;
  wire tie_low_T32Y65;
  wire tie_high_T32Y65;
  wire tie_low_T33Y65;
  wire tie_high_T33Y65;
  wire tie_low_T34Y65;
  wire tie_high_T34Y65;
  wire tie_low_T35Y65;
  wire tie_high_T35Y65;
  wire tie_low_T0Y66;
  wire tie_high_T0Y66;
  wire tie_low_T1Y66;
  wire tie_high_T1Y66;
  wire tie_low_T2Y66;
  wire tie_high_T2Y66;
  wire tie_low_T3Y66;
  wire tie_high_T3Y66;
  wire tie_low_T4Y66;
  wire tie_high_T4Y66;
  wire tie_low_T5Y66;
  wire tie_high_T5Y66;
  wire tie_low_T6Y66;
  wire tie_high_T6Y66;
  wire tie_low_T7Y66;
  wire tie_high_T7Y66;
  wire tie_low_T8Y66;
  wire tie_high_T8Y66;
  wire tie_low_T9Y66;
  wire tie_high_T9Y66;
  wire tie_low_T10Y66;
  wire tie_high_T10Y66;
  wire tie_low_T11Y66;
  wire tie_high_T11Y66;
  wire tie_low_T12Y66;
  wire tie_high_T12Y66;
  wire tie_low_T13Y66;
  wire tie_high_T13Y66;
  wire tie_low_T14Y66;
  wire tie_high_T14Y66;
  wire tie_low_T15Y66;
  wire tie_high_T15Y66;
  wire tie_low_T16Y66;
  wire tie_high_T16Y66;
  wire tie_low_T17Y66;
  wire tie_high_T17Y66;
  wire tie_low_T18Y66;
  wire tie_high_T18Y66;
  wire tie_low_T19Y66;
  wire tie_high_T19Y66;
  wire tie_low_T20Y66;
  wire tie_high_T20Y66;
  wire tie_low_T21Y66;
  wire tie_high_T21Y66;
  wire tie_low_T22Y66;
  wire tie_high_T22Y66;
  wire tie_low_T23Y66;
  wire tie_high_T23Y66;
  wire tie_low_T24Y66;
  wire tie_high_T24Y66;
  wire tie_low_T25Y66;
  wire tie_high_T25Y66;
  wire tie_low_T26Y66;
  wire tie_high_T26Y66;
  wire tie_low_T27Y66;
  wire tie_high_T27Y66;
  wire tie_low_T28Y66;
  wire tie_high_T28Y66;
  wire tie_low_T29Y66;
  wire tie_high_T29Y66;
  wire tie_low_T30Y66;
  wire tie_high_T30Y66;
  wire tie_low_T31Y66;
  wire tie_high_T31Y66;
  wire tie_low_T32Y66;
  wire tie_high_T32Y66;
  wire tie_low_T33Y66;
  wire tie_high_T33Y66;
  wire tie_low_T34Y66;
  wire tie_high_T34Y66;
  wire tie_low_T35Y66;
  wire tie_high_T35Y66;
  wire tie_low_T0Y67;
  wire tie_high_T0Y67;
  wire tie_low_T1Y67;
  wire tie_high_T1Y67;
  wire tie_low_T2Y67;
  wire tie_high_T2Y67;
  wire tie_low_T3Y67;
  wire tie_high_T3Y67;
  wire tie_low_T4Y67;
  wire tie_high_T4Y67;
  wire tie_low_T5Y67;
  wire tie_high_T5Y67;
  wire tie_low_T6Y67;
  wire tie_high_T6Y67;
  wire tie_low_T7Y67;
  wire tie_high_T7Y67;
  wire tie_low_T8Y67;
  wire tie_high_T8Y67;
  wire tie_low_T9Y67;
  wire tie_high_T9Y67;
  wire tie_low_T10Y67;
  wire tie_high_T10Y67;
  wire tie_low_T11Y67;
  wire tie_high_T11Y67;
  wire tie_low_T12Y67;
  wire tie_high_T12Y67;
  wire tie_low_T13Y67;
  wire tie_high_T13Y67;
  wire tie_low_T14Y67;
  wire tie_high_T14Y67;
  wire tie_low_T15Y67;
  wire tie_high_T15Y67;
  wire tie_low_T16Y67;
  wire tie_high_T16Y67;
  wire tie_low_T17Y67;
  wire tie_high_T17Y67;
  wire tie_low_T18Y67;
  wire tie_high_T18Y67;
  wire tie_low_T19Y67;
  wire tie_high_T19Y67;
  wire tie_low_T20Y67;
  wire tie_high_T20Y67;
  wire tie_low_T21Y67;
  wire tie_high_T21Y67;
  wire tie_low_T22Y67;
  wire tie_high_T22Y67;
  wire tie_low_T23Y67;
  wire tie_high_T23Y67;
  wire tie_low_T24Y67;
  wire tie_high_T24Y67;
  wire tie_low_T25Y67;
  wire tie_high_T25Y67;
  wire tie_low_T26Y67;
  wire tie_high_T26Y67;
  wire tie_low_T27Y67;
  wire tie_high_T27Y67;
  wire tie_low_T28Y67;
  wire tie_high_T28Y67;
  wire tie_low_T29Y67;
  wire tie_high_T29Y67;
  wire tie_low_T30Y67;
  wire tie_high_T30Y67;
  wire tie_low_T31Y67;
  wire tie_high_T31Y67;
  wire tie_low_T32Y67;
  wire tie_high_T32Y67;
  wire tie_low_T33Y67;
  wire tie_high_T33Y67;
  wire tie_low_T34Y67;
  wire tie_high_T34Y67;
  wire tie_low_T35Y67;
  wire tie_high_T35Y67;
  wire tie_low_T0Y68;
  wire tie_high_T0Y68;
  wire tie_low_T1Y68;
  wire tie_high_T1Y68;
  wire tie_low_T2Y68;
  wire tie_high_T2Y68;
  wire tie_low_T3Y68;
  wire tie_high_T3Y68;
  wire tie_low_T4Y68;
  wire tie_high_T4Y68;
  wire tie_low_T5Y68;
  wire tie_high_T5Y68;
  wire tie_low_T6Y68;
  wire tie_high_T6Y68;
  wire tie_low_T7Y68;
  wire tie_high_T7Y68;
  wire tie_low_T8Y68;
  wire tie_high_T8Y68;
  wire tie_low_T9Y68;
  wire tie_high_T9Y68;
  wire tie_low_T10Y68;
  wire tie_high_T10Y68;
  wire tie_low_T11Y68;
  wire tie_high_T11Y68;
  wire tie_low_T12Y68;
  wire tie_high_T12Y68;
  wire tie_low_T13Y68;
  wire tie_high_T13Y68;
  wire tie_low_T14Y68;
  wire tie_high_T14Y68;
  wire tie_low_T15Y68;
  wire tie_high_T15Y68;
  wire tie_low_T16Y68;
  wire tie_high_T16Y68;
  wire tie_low_T17Y68;
  wire tie_high_T17Y68;
  wire tie_low_T18Y68;
  wire tie_high_T18Y68;
  wire tie_low_T19Y68;
  wire tie_high_T19Y68;
  wire tie_low_T20Y68;
  wire tie_high_T20Y68;
  wire tie_low_T21Y68;
  wire tie_high_T21Y68;
  wire tie_low_T22Y68;
  wire tie_high_T22Y68;
  wire tie_low_T23Y68;
  wire tie_high_T23Y68;
  wire tie_low_T24Y68;
  wire tie_high_T24Y68;
  wire tie_low_T25Y68;
  wire tie_high_T25Y68;
  wire tie_low_T26Y68;
  wire tie_high_T26Y68;
  wire tie_low_T27Y68;
  wire tie_high_T27Y68;
  wire tie_low_T28Y68;
  wire tie_high_T28Y68;
  wire tie_low_T29Y68;
  wire tie_high_T29Y68;
  wire tie_low_T30Y68;
  wire tie_high_T30Y68;
  wire tie_low_T31Y68;
  wire tie_high_T31Y68;
  wire tie_low_T32Y68;
  wire tie_high_T32Y68;
  wire tie_low_T33Y68;
  wire tie_high_T33Y68;
  wire tie_low_T34Y68;
  wire tie_high_T34Y68;
  wire tie_low_T35Y68;
  wire tie_high_T35Y68;
  wire tie_low_T0Y69;
  wire tie_high_T0Y69;
  wire tie_low_T1Y69;
  wire tie_high_T1Y69;
  wire tie_low_T2Y69;
  wire tie_high_T2Y69;
  wire tie_low_T3Y69;
  wire tie_high_T3Y69;
  wire tie_low_T4Y69;
  wire tie_high_T4Y69;
  wire tie_low_T5Y69;
  wire tie_high_T5Y69;
  wire tie_low_T6Y69;
  wire tie_high_T6Y69;
  wire tie_low_T7Y69;
  wire tie_high_T7Y69;
  wire tie_low_T8Y69;
  wire tie_high_T8Y69;
  wire tie_low_T9Y69;
  wire tie_high_T9Y69;
  wire tie_low_T10Y69;
  wire tie_high_T10Y69;
  wire tie_low_T11Y69;
  wire tie_high_T11Y69;
  wire tie_low_T12Y69;
  wire tie_high_T12Y69;
  wire tie_low_T13Y69;
  wire tie_high_T13Y69;
  wire tie_low_T14Y69;
  wire tie_high_T14Y69;
  wire tie_low_T15Y69;
  wire tie_high_T15Y69;
  wire tie_low_T16Y69;
  wire tie_high_T16Y69;
  wire tie_low_T17Y69;
  wire tie_high_T17Y69;
  wire tie_low_T18Y69;
  wire tie_high_T18Y69;
  wire tie_low_T19Y69;
  wire tie_high_T19Y69;
  wire tie_low_T20Y69;
  wire tie_high_T20Y69;
  wire tie_low_T21Y69;
  wire tie_high_T21Y69;
  wire tie_low_T22Y69;
  wire tie_high_T22Y69;
  wire tie_low_T23Y69;
  wire tie_high_T23Y69;
  wire tie_low_T24Y69;
  wire tie_high_T24Y69;
  wire tie_low_T25Y69;
  wire tie_high_T25Y69;
  wire tie_low_T26Y69;
  wire tie_high_T26Y69;
  wire tie_low_T27Y69;
  wire tie_high_T27Y69;
  wire tie_low_T28Y69;
  wire tie_high_T28Y69;
  wire tie_low_T29Y69;
  wire tie_high_T29Y69;
  wire tie_low_T30Y69;
  wire tie_high_T30Y69;
  wire tie_low_T31Y69;
  wire tie_high_T31Y69;
  wire tie_low_T32Y69;
  wire tie_high_T32Y69;
  wire tie_low_T33Y69;
  wire tie_high_T33Y69;
  wire tie_low_T34Y69;
  wire tie_high_T34Y69;
  wire tie_low_T35Y69;
  wire tie_high_T35Y69;
  wire tie_low_T0Y70;
  wire tie_high_T0Y70;
  wire tie_low_T1Y70;
  wire tie_high_T1Y70;
  wire tie_low_T2Y70;
  wire tie_high_T2Y70;
  wire tie_low_T3Y70;
  wire tie_high_T3Y70;
  wire tie_low_T4Y70;
  wire tie_high_T4Y70;
  wire tie_low_T5Y70;
  wire tie_high_T5Y70;
  wire tie_low_T6Y70;
  wire tie_high_T6Y70;
  wire tie_low_T7Y70;
  wire tie_high_T7Y70;
  wire tie_low_T8Y70;
  wire tie_high_T8Y70;
  wire tie_low_T9Y70;
  wire tie_high_T9Y70;
  wire tie_low_T10Y70;
  wire tie_high_T10Y70;
  wire tie_low_T11Y70;
  wire tie_high_T11Y70;
  wire tie_low_T12Y70;
  wire tie_high_T12Y70;
  wire tie_low_T13Y70;
  wire tie_high_T13Y70;
  wire tie_low_T14Y70;
  wire tie_high_T14Y70;
  wire tie_low_T15Y70;
  wire tie_high_T15Y70;
  wire tie_low_T16Y70;
  wire tie_high_T16Y70;
  wire tie_low_T17Y70;
  wire tie_high_T17Y70;
  wire tie_low_T18Y70;
  wire tie_high_T18Y70;
  wire tie_low_T19Y70;
  wire tie_high_T19Y70;
  wire tie_low_T20Y70;
  wire tie_high_T20Y70;
  wire tie_low_T21Y70;
  wire tie_high_T21Y70;
  wire tie_low_T22Y70;
  wire tie_high_T22Y70;
  wire tie_low_T23Y70;
  wire tie_high_T23Y70;
  wire tie_low_T24Y70;
  wire tie_high_T24Y70;
  wire tie_low_T25Y70;
  wire tie_high_T25Y70;
  wire tie_low_T26Y70;
  wire tie_high_T26Y70;
  wire tie_low_T27Y70;
  wire tie_high_T27Y70;
  wire tie_low_T28Y70;
  wire tie_high_T28Y70;
  wire tie_low_T29Y70;
  wire tie_high_T29Y70;
  wire tie_low_T30Y70;
  wire tie_high_T30Y70;
  wire tie_low_T31Y70;
  wire tie_high_T31Y70;
  wire tie_low_T32Y70;
  wire tie_high_T32Y70;
  wire tie_low_T33Y70;
  wire tie_high_T33Y70;
  wire tie_low_T34Y70;
  wire tie_high_T34Y70;
  wire tie_low_T35Y70;
  wire tie_high_T35Y70;
  wire tie_low_T0Y71;
  wire tie_high_T0Y71;
  wire tie_low_T1Y71;
  wire tie_high_T1Y71;
  wire tie_low_T2Y71;
  wire tie_high_T2Y71;
  wire tie_low_T3Y71;
  wire tie_high_T3Y71;
  wire tie_low_T4Y71;
  wire tie_high_T4Y71;
  wire tie_low_T5Y71;
  wire tie_high_T5Y71;
  wire tie_low_T6Y71;
  wire tie_high_T6Y71;
  wire tie_low_T7Y71;
  wire tie_high_T7Y71;
  wire tie_low_T8Y71;
  wire tie_high_T8Y71;
  wire tie_low_T9Y71;
  wire tie_high_T9Y71;
  wire tie_low_T10Y71;
  wire tie_high_T10Y71;
  wire tie_low_T11Y71;
  wire tie_high_T11Y71;
  wire tie_low_T12Y71;
  wire tie_high_T12Y71;
  wire tie_low_T13Y71;
  wire tie_high_T13Y71;
  wire tie_low_T14Y71;
  wire tie_high_T14Y71;
  wire tie_low_T15Y71;
  wire tie_high_T15Y71;
  wire tie_low_T16Y71;
  wire tie_high_T16Y71;
  wire tie_low_T17Y71;
  wire tie_high_T17Y71;
  wire tie_low_T18Y71;
  wire tie_high_T18Y71;
  wire tie_low_T19Y71;
  wire tie_high_T19Y71;
  wire tie_low_T20Y71;
  wire tie_high_T20Y71;
  wire tie_low_T21Y71;
  wire tie_high_T21Y71;
  wire tie_low_T22Y71;
  wire tie_high_T22Y71;
  wire tie_low_T23Y71;
  wire tie_high_T23Y71;
  wire tie_low_T24Y71;
  wire tie_high_T24Y71;
  wire tie_low_T25Y71;
  wire tie_high_T25Y71;
  wire tie_low_T26Y71;
  wire tie_high_T26Y71;
  wire tie_low_T27Y71;
  wire tie_high_T27Y71;
  wire tie_low_T28Y71;
  wire tie_high_T28Y71;
  wire tie_low_T29Y71;
  wire tie_high_T29Y71;
  wire tie_low_T30Y71;
  wire tie_high_T30Y71;
  wire tie_low_T31Y71;
  wire tie_high_T31Y71;
  wire tie_low_T32Y71;
  wire tie_high_T32Y71;
  wire tie_low_T33Y71;
  wire tie_high_T33Y71;
  wire tie_low_T34Y71;
  wire tie_high_T34Y71;
  wire tie_low_T35Y71;
  wire tie_high_T35Y71;
  wire tie_low_T0Y72;
  wire tie_high_T0Y72;
  wire tie_low_T1Y72;
  wire tie_high_T1Y72;
  wire tie_low_T2Y72;
  wire tie_high_T2Y72;
  wire tie_low_T3Y72;
  wire tie_high_T3Y72;
  wire tie_low_T4Y72;
  wire tie_high_T4Y72;
  wire tie_low_T5Y72;
  wire tie_high_T5Y72;
  wire tie_low_T6Y72;
  wire tie_high_T6Y72;
  wire tie_low_T7Y72;
  wire tie_high_T7Y72;
  wire tie_low_T8Y72;
  wire tie_high_T8Y72;
  wire tie_low_T9Y72;
  wire tie_high_T9Y72;
  wire tie_low_T10Y72;
  wire tie_high_T10Y72;
  wire tie_low_T11Y72;
  wire tie_high_T11Y72;
  wire tie_low_T12Y72;
  wire tie_high_T12Y72;
  wire tie_low_T13Y72;
  wire tie_high_T13Y72;
  wire tie_low_T14Y72;
  wire tie_high_T14Y72;
  wire tie_low_T15Y72;
  wire tie_high_T15Y72;
  wire tie_low_T16Y72;
  wire tie_high_T16Y72;
  wire tie_low_T17Y72;
  wire tie_high_T17Y72;
  wire tie_low_T18Y72;
  wire tie_high_T18Y72;
  wire tie_low_T19Y72;
  wire tie_high_T19Y72;
  wire tie_low_T20Y72;
  wire tie_high_T20Y72;
  wire tie_low_T21Y72;
  wire tie_high_T21Y72;
  wire tie_low_T22Y72;
  wire tie_high_T22Y72;
  wire tie_low_T23Y72;
  wire tie_high_T23Y72;
  wire tie_low_T24Y72;
  wire tie_high_T24Y72;
  wire tie_low_T25Y72;
  wire tie_high_T25Y72;
  wire tie_low_T26Y72;
  wire tie_high_T26Y72;
  wire tie_low_T27Y72;
  wire tie_high_T27Y72;
  wire tie_low_T28Y72;
  wire tie_high_T28Y72;
  wire tie_low_T29Y72;
  wire tie_high_T29Y72;
  wire tie_low_T30Y72;
  wire tie_high_T30Y72;
  wire tie_low_T31Y72;
  wire tie_high_T31Y72;
  wire tie_low_T32Y72;
  wire tie_high_T32Y72;
  wire tie_low_T33Y72;
  wire tie_high_T33Y72;
  wire tie_low_T34Y72;
  wire tie_high_T34Y72;
  wire tie_low_T35Y72;
  wire tie_high_T35Y72;
  wire tie_low_T0Y73;
  wire tie_high_T0Y73;
  wire tie_low_T1Y73;
  wire tie_high_T1Y73;
  wire tie_low_T2Y73;
  wire tie_high_T2Y73;
  wire tie_low_T3Y73;
  wire tie_high_T3Y73;
  wire tie_low_T4Y73;
  wire tie_high_T4Y73;
  wire tie_low_T5Y73;
  wire tie_high_T5Y73;
  wire tie_low_T6Y73;
  wire tie_high_T6Y73;
  wire tie_low_T7Y73;
  wire tie_high_T7Y73;
  wire tie_low_T8Y73;
  wire tie_high_T8Y73;
  wire tie_low_T9Y73;
  wire tie_high_T9Y73;
  wire tie_low_T10Y73;
  wire tie_high_T10Y73;
  wire tie_low_T11Y73;
  wire tie_high_T11Y73;
  wire tie_low_T12Y73;
  wire tie_high_T12Y73;
  wire tie_low_T13Y73;
  wire tie_high_T13Y73;
  wire tie_low_T14Y73;
  wire tie_high_T14Y73;
  wire tie_low_T15Y73;
  wire tie_high_T15Y73;
  wire tie_low_T16Y73;
  wire tie_high_T16Y73;
  wire tie_low_T17Y73;
  wire tie_high_T17Y73;
  wire tie_low_T18Y73;
  wire tie_high_T18Y73;
  wire tie_low_T19Y73;
  wire tie_high_T19Y73;
  wire tie_low_T20Y73;
  wire tie_high_T20Y73;
  wire tie_low_T21Y73;
  wire tie_high_T21Y73;
  wire tie_low_T22Y73;
  wire tie_high_T22Y73;
  wire tie_low_T23Y73;
  wire tie_high_T23Y73;
  wire tie_low_T24Y73;
  wire tie_high_T24Y73;
  wire tie_low_T25Y73;
  wire tie_high_T25Y73;
  wire tie_low_T26Y73;
  wire tie_high_T26Y73;
  wire tie_low_T27Y73;
  wire tie_high_T27Y73;
  wire tie_low_T28Y73;
  wire tie_high_T28Y73;
  wire tie_low_T29Y73;
  wire tie_high_T29Y73;
  wire tie_low_T30Y73;
  wire tie_high_T30Y73;
  wire tie_low_T31Y73;
  wire tie_high_T31Y73;
  wire tie_low_T32Y73;
  wire tie_high_T32Y73;
  wire tie_low_T33Y73;
  wire tie_high_T33Y73;
  wire tie_low_T34Y73;
  wire tie_high_T34Y73;
  wire tie_low_T35Y73;
  wire tie_high_T35Y73;
  wire tie_low_T0Y74;
  wire tie_high_T0Y74;
  wire tie_low_T1Y74;
  wire tie_high_T1Y74;
  wire tie_low_T2Y74;
  wire tie_high_T2Y74;
  wire tie_low_T3Y74;
  wire tie_high_T3Y74;
  wire tie_low_T4Y74;
  wire tie_high_T4Y74;
  wire tie_low_T5Y74;
  wire tie_high_T5Y74;
  wire tie_low_T6Y74;
  wire tie_high_T6Y74;
  wire tie_low_T7Y74;
  wire tie_high_T7Y74;
  wire tie_low_T8Y74;
  wire tie_high_T8Y74;
  wire tie_low_T9Y74;
  wire tie_high_T9Y74;
  wire tie_low_T10Y74;
  wire tie_high_T10Y74;
  wire tie_low_T11Y74;
  wire tie_high_T11Y74;
  wire tie_low_T12Y74;
  wire tie_high_T12Y74;
  wire tie_low_T13Y74;
  wire tie_high_T13Y74;
  wire tie_low_T14Y74;
  wire tie_high_T14Y74;
  wire tie_low_T15Y74;
  wire tie_high_T15Y74;
  wire tie_low_T16Y74;
  wire tie_high_T16Y74;
  wire tie_low_T17Y74;
  wire tie_high_T17Y74;
  wire tie_low_T18Y74;
  wire tie_high_T18Y74;
  wire tie_low_T19Y74;
  wire tie_high_T19Y74;
  wire tie_low_T20Y74;
  wire tie_high_T20Y74;
  wire tie_low_T21Y74;
  wire tie_high_T21Y74;
  wire tie_low_T22Y74;
  wire tie_high_T22Y74;
  wire tie_low_T23Y74;
  wire tie_high_T23Y74;
  wire tie_low_T24Y74;
  wire tie_high_T24Y74;
  wire tie_low_T25Y74;
  wire tie_high_T25Y74;
  wire tie_low_T26Y74;
  wire tie_high_T26Y74;
  wire tie_low_T27Y74;
  wire tie_high_T27Y74;
  wire tie_low_T28Y74;
  wire tie_high_T28Y74;
  wire tie_low_T29Y74;
  wire tie_high_T29Y74;
  wire tie_low_T30Y74;
  wire tie_high_T30Y74;
  wire tie_low_T31Y74;
  wire tie_high_T31Y74;
  wire tie_low_T32Y74;
  wire tie_high_T32Y74;
  wire tie_low_T33Y74;
  wire tie_high_T33Y74;
  wire tie_low_T34Y74;
  wire tie_high_T34Y74;
  wire tie_low_T35Y74;
  wire tie_high_T35Y74;
  wire tie_low_T0Y75;
  wire tie_high_T0Y75;
  wire tie_low_T1Y75;
  wire tie_high_T1Y75;
  wire tie_low_T2Y75;
  wire tie_high_T2Y75;
  wire tie_low_T3Y75;
  wire tie_high_T3Y75;
  wire tie_low_T4Y75;
  wire tie_high_T4Y75;
  wire tie_low_T5Y75;
  wire tie_high_T5Y75;
  wire tie_low_T6Y75;
  wire tie_high_T6Y75;
  wire tie_low_T7Y75;
  wire tie_high_T7Y75;
  wire tie_low_T8Y75;
  wire tie_high_T8Y75;
  wire tie_low_T9Y75;
  wire tie_high_T9Y75;
  wire tie_low_T10Y75;
  wire tie_high_T10Y75;
  wire tie_low_T11Y75;
  wire tie_high_T11Y75;
  wire tie_low_T12Y75;
  wire tie_high_T12Y75;
  wire tie_low_T13Y75;
  wire tie_high_T13Y75;
  wire tie_low_T14Y75;
  wire tie_high_T14Y75;
  wire tie_low_T15Y75;
  wire tie_high_T15Y75;
  wire tie_low_T16Y75;
  wire tie_high_T16Y75;
  wire tie_low_T17Y75;
  wire tie_high_T17Y75;
  wire tie_low_T18Y75;
  wire tie_high_T18Y75;
  wire tie_low_T19Y75;
  wire tie_high_T19Y75;
  wire tie_low_T20Y75;
  wire tie_high_T20Y75;
  wire tie_low_T21Y75;
  wire tie_high_T21Y75;
  wire tie_low_T22Y75;
  wire tie_high_T22Y75;
  wire tie_low_T23Y75;
  wire tie_high_T23Y75;
  wire tie_low_T24Y75;
  wire tie_high_T24Y75;
  wire tie_low_T25Y75;
  wire tie_high_T25Y75;
  wire tie_low_T26Y75;
  wire tie_high_T26Y75;
  wire tie_low_T27Y75;
  wire tie_high_T27Y75;
  wire tie_low_T28Y75;
  wire tie_high_T28Y75;
  wire tie_low_T29Y75;
  wire tie_high_T29Y75;
  wire tie_low_T30Y75;
  wire tie_high_T30Y75;
  wire tie_low_T31Y75;
  wire tie_high_T31Y75;
  wire tie_low_T32Y75;
  wire tie_high_T32Y75;
  wire tie_low_T33Y75;
  wire tie_high_T33Y75;
  wire tie_low_T34Y75;
  wire tie_high_T34Y75;
  wire tie_low_T35Y75;
  wire tie_high_T35Y75;
  wire tie_low_T0Y76;
  wire tie_high_T0Y76;
  wire tie_low_T1Y76;
  wire tie_high_T1Y76;
  wire tie_low_T2Y76;
  wire tie_high_T2Y76;
  wire tie_low_T3Y76;
  wire tie_high_T3Y76;
  wire tie_low_T4Y76;
  wire tie_high_T4Y76;
  wire tie_low_T5Y76;
  wire tie_high_T5Y76;
  wire tie_low_T6Y76;
  wire tie_high_T6Y76;
  wire tie_low_T7Y76;
  wire tie_high_T7Y76;
  wire tie_low_T8Y76;
  wire tie_high_T8Y76;
  wire tie_low_T9Y76;
  wire tie_high_T9Y76;
  wire tie_low_T10Y76;
  wire tie_high_T10Y76;
  wire tie_low_T11Y76;
  wire tie_high_T11Y76;
  wire tie_low_T12Y76;
  wire tie_high_T12Y76;
  wire tie_low_T13Y76;
  wire tie_high_T13Y76;
  wire tie_low_T14Y76;
  wire tie_high_T14Y76;
  wire tie_low_T15Y76;
  wire tie_high_T15Y76;
  wire tie_low_T16Y76;
  wire tie_high_T16Y76;
  wire tie_low_T17Y76;
  wire tie_high_T17Y76;
  wire tie_low_T18Y76;
  wire tie_high_T18Y76;
  wire tie_low_T19Y76;
  wire tie_high_T19Y76;
  wire tie_low_T20Y76;
  wire tie_high_T20Y76;
  wire tie_low_T21Y76;
  wire tie_high_T21Y76;
  wire tie_low_T22Y76;
  wire tie_high_T22Y76;
  wire tie_low_T23Y76;
  wire tie_high_T23Y76;
  wire tie_low_T24Y76;
  wire tie_high_T24Y76;
  wire tie_low_T25Y76;
  wire tie_high_T25Y76;
  wire tie_low_T26Y76;
  wire tie_high_T26Y76;
  wire tie_low_T27Y76;
  wire tie_high_T27Y76;
  wire tie_low_T28Y76;
  wire tie_high_T28Y76;
  wire tie_low_T29Y76;
  wire tie_high_T29Y76;
  wire tie_low_T30Y76;
  wire tie_high_T30Y76;
  wire tie_low_T31Y76;
  wire tie_high_T31Y76;
  wire tie_low_T32Y76;
  wire tie_high_T32Y76;
  wire tie_low_T33Y76;
  wire tie_high_T33Y76;
  wire tie_low_T34Y76;
  wire tie_high_T34Y76;
  wire tie_low_T35Y76;
  wire tie_high_T35Y76;
  wire tie_low_T0Y77;
  wire tie_high_T0Y77;
  wire tie_low_T1Y77;
  wire tie_high_T1Y77;
  wire tie_low_T2Y77;
  wire tie_high_T2Y77;
  wire tie_low_T3Y77;
  wire tie_high_T3Y77;
  wire tie_low_T4Y77;
  wire tie_high_T4Y77;
  wire tie_low_T5Y77;
  wire tie_high_T5Y77;
  wire tie_low_T6Y77;
  wire tie_high_T6Y77;
  wire tie_low_T7Y77;
  wire tie_high_T7Y77;
  wire tie_low_T8Y77;
  wire tie_high_T8Y77;
  wire tie_low_T9Y77;
  wire tie_high_T9Y77;
  wire tie_low_T10Y77;
  wire tie_high_T10Y77;
  wire tie_low_T11Y77;
  wire tie_high_T11Y77;
  wire tie_low_T12Y77;
  wire tie_high_T12Y77;
  wire tie_low_T13Y77;
  wire tie_high_T13Y77;
  wire tie_low_T14Y77;
  wire tie_high_T14Y77;
  wire tie_low_T15Y77;
  wire tie_high_T15Y77;
  wire tie_low_T16Y77;
  wire tie_high_T16Y77;
  wire tie_low_T17Y77;
  wire tie_high_T17Y77;
  wire tie_low_T18Y77;
  wire tie_high_T18Y77;
  wire tie_low_T19Y77;
  wire tie_high_T19Y77;
  wire tie_low_T20Y77;
  wire tie_high_T20Y77;
  wire tie_low_T21Y77;
  wire tie_high_T21Y77;
  wire tie_low_T22Y77;
  wire tie_high_T22Y77;
  wire tie_low_T23Y77;
  wire tie_high_T23Y77;
  wire tie_low_T24Y77;
  wire tie_high_T24Y77;
  wire tie_low_T25Y77;
  wire tie_high_T25Y77;
  wire tie_low_T26Y77;
  wire tie_high_T26Y77;
  wire tie_low_T27Y77;
  wire tie_high_T27Y77;
  wire tie_low_T28Y77;
  wire tie_high_T28Y77;
  wire tie_low_T29Y77;
  wire tie_high_T29Y77;
  wire tie_low_T30Y77;
  wire tie_high_T30Y77;
  wire tie_low_T31Y77;
  wire tie_high_T31Y77;
  wire tie_low_T32Y77;
  wire tie_high_T32Y77;
  wire tie_low_T33Y77;
  wire tie_high_T33Y77;
  wire tie_low_T34Y77;
  wire tie_high_T34Y77;
  wire tie_low_T35Y77;
  wire tie_high_T35Y77;
  wire tie_low_T0Y78;
  wire tie_high_T0Y78;
  wire tie_low_T1Y78;
  wire tie_high_T1Y78;
  wire tie_low_T2Y78;
  wire tie_high_T2Y78;
  wire tie_low_T3Y78;
  wire tie_high_T3Y78;
  wire tie_low_T4Y78;
  wire tie_high_T4Y78;
  wire tie_low_T5Y78;
  wire tie_high_T5Y78;
  wire tie_low_T6Y78;
  wire tie_high_T6Y78;
  wire tie_low_T7Y78;
  wire tie_high_T7Y78;
  wire tie_low_T8Y78;
  wire tie_high_T8Y78;
  wire tie_low_T9Y78;
  wire tie_high_T9Y78;
  wire tie_low_T10Y78;
  wire tie_high_T10Y78;
  wire tie_low_T11Y78;
  wire tie_high_T11Y78;
  wire tie_low_T12Y78;
  wire tie_high_T12Y78;
  wire tie_low_T13Y78;
  wire tie_high_T13Y78;
  wire tie_low_T14Y78;
  wire tie_high_T14Y78;
  wire tie_low_T15Y78;
  wire tie_high_T15Y78;
  wire tie_low_T16Y78;
  wire tie_high_T16Y78;
  wire tie_low_T17Y78;
  wire tie_high_T17Y78;
  wire tie_low_T18Y78;
  wire tie_high_T18Y78;
  wire tie_low_T19Y78;
  wire tie_high_T19Y78;
  wire tie_low_T20Y78;
  wire tie_high_T20Y78;
  wire tie_low_T21Y78;
  wire tie_high_T21Y78;
  wire tie_low_T22Y78;
  wire tie_high_T22Y78;
  wire tie_low_T23Y78;
  wire tie_high_T23Y78;
  wire tie_low_T24Y78;
  wire tie_high_T24Y78;
  wire tie_low_T25Y78;
  wire tie_high_T25Y78;
  wire tie_low_T26Y78;
  wire tie_high_T26Y78;
  wire tie_low_T27Y78;
  wire tie_high_T27Y78;
  wire tie_low_T28Y78;
  wire tie_high_T28Y78;
  wire tie_low_T29Y78;
  wire tie_high_T29Y78;
  wire tie_low_T30Y78;
  wire tie_high_T30Y78;
  wire tie_low_T31Y78;
  wire tie_high_T31Y78;
  wire tie_low_T32Y78;
  wire tie_high_T32Y78;
  wire tie_low_T33Y78;
  wire tie_high_T33Y78;
  wire tie_low_T34Y78;
  wire tie_high_T34Y78;
  wire tie_low_T35Y78;
  wire tie_high_T35Y78;
  wire tie_low_T0Y79;
  wire tie_high_T0Y79;
  wire tie_low_T1Y79;
  wire tie_high_T1Y79;
  wire tie_low_T2Y79;
  wire tie_high_T2Y79;
  wire tie_low_T3Y79;
  wire tie_high_T3Y79;
  wire tie_low_T4Y79;
  wire tie_high_T4Y79;
  wire tie_low_T5Y79;
  wire tie_high_T5Y79;
  wire tie_low_T6Y79;
  wire tie_high_T6Y79;
  wire tie_low_T7Y79;
  wire tie_high_T7Y79;
  wire tie_low_T8Y79;
  wire tie_high_T8Y79;
  wire tie_low_T9Y79;
  wire tie_high_T9Y79;
  wire tie_low_T10Y79;
  wire tie_high_T10Y79;
  wire tie_low_T11Y79;
  wire tie_high_T11Y79;
  wire tie_low_T12Y79;
  wire tie_high_T12Y79;
  wire tie_low_T13Y79;
  wire tie_high_T13Y79;
  wire tie_low_T14Y79;
  wire tie_high_T14Y79;
  wire tie_low_T15Y79;
  wire tie_high_T15Y79;
  wire tie_low_T16Y79;
  wire tie_high_T16Y79;
  wire tie_low_T17Y79;
  wire tie_high_T17Y79;
  wire tie_low_T18Y79;
  wire tie_high_T18Y79;
  wire tie_low_T19Y79;
  wire tie_high_T19Y79;
  wire tie_low_T20Y79;
  wire tie_high_T20Y79;
  wire tie_low_T21Y79;
  wire tie_high_T21Y79;
  wire tie_low_T22Y79;
  wire tie_high_T22Y79;
  wire tie_low_T23Y79;
  wire tie_high_T23Y79;
  wire tie_low_T24Y79;
  wire tie_high_T24Y79;
  wire tie_low_T25Y79;
  wire tie_high_T25Y79;
  wire tie_low_T26Y79;
  wire tie_high_T26Y79;
  wire tie_low_T27Y79;
  wire tie_high_T27Y79;
  wire tie_low_T28Y79;
  wire tie_high_T28Y79;
  wire tie_low_T29Y79;
  wire tie_high_T29Y79;
  wire tie_low_T30Y79;
  wire tie_high_T30Y79;
  wire tie_low_T31Y79;
  wire tie_high_T31Y79;
  wire tie_low_T32Y79;
  wire tie_high_T32Y79;
  wire tie_low_T33Y79;
  wire tie_high_T33Y79;
  wire tie_low_T34Y79;
  wire tie_high_T34Y79;
  wire tie_low_T35Y79;
  wire tie_high_T35Y79;
  wire tie_low_T0Y80;
  wire tie_high_T0Y80;
  wire tie_low_T1Y80;
  wire tie_high_T1Y80;
  wire tie_low_T2Y80;
  wire tie_high_T2Y80;
  wire tie_low_T3Y80;
  wire tie_high_T3Y80;
  wire tie_low_T4Y80;
  wire tie_high_T4Y80;
  wire tie_low_T5Y80;
  wire tie_high_T5Y80;
  wire tie_low_T6Y80;
  wire tie_high_T6Y80;
  wire tie_low_T7Y80;
  wire tie_high_T7Y80;
  wire tie_low_T8Y80;
  wire tie_high_T8Y80;
  wire tie_low_T9Y80;
  wire tie_high_T9Y80;
  wire tie_low_T10Y80;
  wire tie_high_T10Y80;
  wire tie_low_T11Y80;
  wire tie_high_T11Y80;
  wire tie_low_T12Y80;
  wire tie_high_T12Y80;
  wire tie_low_T13Y80;
  wire tie_high_T13Y80;
  wire tie_low_T14Y80;
  wire tie_high_T14Y80;
  wire tie_low_T15Y80;
  wire tie_high_T15Y80;
  wire tie_low_T16Y80;
  wire tie_high_T16Y80;
  wire tie_low_T17Y80;
  wire tie_high_T17Y80;
  wire tie_low_T18Y80;
  wire tie_high_T18Y80;
  wire tie_low_T19Y80;
  wire tie_high_T19Y80;
  wire tie_low_T20Y80;
  wire tie_high_T20Y80;
  wire tie_low_T21Y80;
  wire tie_high_T21Y80;
  wire tie_low_T22Y80;
  wire tie_high_T22Y80;
  wire tie_low_T23Y80;
  wire tie_high_T23Y80;
  wire tie_low_T24Y80;
  wire tie_high_T24Y80;
  wire tie_low_T25Y80;
  wire tie_high_T25Y80;
  wire tie_low_T26Y80;
  wire tie_high_T26Y80;
  wire tie_low_T27Y80;
  wire tie_high_T27Y80;
  wire tie_low_T28Y80;
  wire tie_high_T28Y80;
  wire tie_low_T29Y80;
  wire tie_high_T29Y80;
  wire tie_low_T30Y80;
  wire tie_high_T30Y80;
  wire tie_low_T31Y80;
  wire tie_high_T31Y80;
  wire tie_low_T32Y80;
  wire tie_high_T32Y80;
  wire tie_low_T33Y80;
  wire tie_high_T33Y80;
  wire tie_low_T34Y80;
  wire tie_high_T34Y80;
  wire tie_low_T35Y80;
  wire tie_high_T35Y80;
  wire tie_low_T0Y81;
  wire tie_high_T0Y81;
  wire tie_low_T1Y81;
  wire tie_high_T1Y81;
  wire tie_low_T2Y81;
  wire tie_high_T2Y81;
  wire tie_low_T3Y81;
  wire tie_high_T3Y81;
  wire tie_low_T4Y81;
  wire tie_high_T4Y81;
  wire tie_low_T5Y81;
  wire tie_high_T5Y81;
  wire tie_low_T6Y81;
  wire tie_high_T6Y81;
  wire tie_low_T7Y81;
  wire tie_high_T7Y81;
  wire tie_low_T8Y81;
  wire tie_high_T8Y81;
  wire tie_low_T9Y81;
  wire tie_high_T9Y81;
  wire tie_low_T10Y81;
  wire tie_high_T10Y81;
  wire tie_low_T11Y81;
  wire tie_high_T11Y81;
  wire tie_low_T12Y81;
  wire tie_high_T12Y81;
  wire tie_low_T13Y81;
  wire tie_high_T13Y81;
  wire tie_low_T14Y81;
  wire tie_high_T14Y81;
  wire tie_low_T15Y81;
  wire tie_high_T15Y81;
  wire tie_low_T16Y81;
  wire tie_high_T16Y81;
  wire tie_low_T17Y81;
  wire tie_high_T17Y81;
  wire tie_low_T18Y81;
  wire tie_high_T18Y81;
  wire tie_low_T19Y81;
  wire tie_high_T19Y81;
  wire tie_low_T20Y81;
  wire tie_high_T20Y81;
  wire tie_low_T21Y81;
  wire tie_high_T21Y81;
  wire tie_low_T22Y81;
  wire tie_high_T22Y81;
  wire tie_low_T23Y81;
  wire tie_high_T23Y81;
  wire tie_low_T24Y81;
  wire tie_high_T24Y81;
  wire tie_low_T25Y81;
  wire tie_high_T25Y81;
  wire tie_low_T26Y81;
  wire tie_high_T26Y81;
  wire tie_low_T27Y81;
  wire tie_high_T27Y81;
  wire tie_low_T28Y81;
  wire tie_high_T28Y81;
  wire tie_low_T29Y81;
  wire tie_high_T29Y81;
  wire tie_low_T30Y81;
  wire tie_high_T30Y81;
  wire tie_low_T31Y81;
  wire tie_high_T31Y81;
  wire tie_low_T32Y81;
  wire tie_high_T32Y81;
  wire tie_low_T33Y81;
  wire tie_high_T33Y81;
  wire tie_low_T34Y81;
  wire tie_high_T34Y81;
  wire tie_low_T35Y81;
  wire tie_high_T35Y81;
  wire tie_low_T0Y82;
  wire tie_high_T0Y82;
  wire tie_low_T1Y82;
  wire tie_high_T1Y82;
  wire tie_low_T2Y82;
  wire tie_high_T2Y82;
  wire tie_low_T3Y82;
  wire tie_high_T3Y82;
  wire tie_low_T4Y82;
  wire tie_high_T4Y82;
  wire tie_low_T5Y82;
  wire tie_high_T5Y82;
  wire tie_low_T6Y82;
  wire tie_high_T6Y82;
  wire tie_low_T7Y82;
  wire tie_high_T7Y82;
  wire tie_low_T8Y82;
  wire tie_high_T8Y82;
  wire tie_low_T9Y82;
  wire tie_high_T9Y82;
  wire tie_low_T10Y82;
  wire tie_high_T10Y82;
  wire tie_low_T11Y82;
  wire tie_high_T11Y82;
  wire tie_low_T12Y82;
  wire tie_high_T12Y82;
  wire tie_low_T13Y82;
  wire tie_high_T13Y82;
  wire tie_low_T14Y82;
  wire tie_high_T14Y82;
  wire tie_low_T15Y82;
  wire tie_high_T15Y82;
  wire tie_low_T16Y82;
  wire tie_high_T16Y82;
  wire tie_low_T17Y82;
  wire tie_high_T17Y82;
  wire tie_low_T18Y82;
  wire tie_high_T18Y82;
  wire tie_low_T19Y82;
  wire tie_high_T19Y82;
  wire tie_low_T20Y82;
  wire tie_high_T20Y82;
  wire tie_low_T21Y82;
  wire tie_high_T21Y82;
  wire tie_low_T22Y82;
  wire tie_high_T22Y82;
  wire tie_low_T23Y82;
  wire tie_high_T23Y82;
  wire tie_low_T24Y82;
  wire tie_high_T24Y82;
  wire tie_low_T25Y82;
  wire tie_high_T25Y82;
  wire tie_low_T26Y82;
  wire tie_high_T26Y82;
  wire tie_low_T27Y82;
  wire tie_high_T27Y82;
  wire tie_low_T28Y82;
  wire tie_high_T28Y82;
  wire tie_low_T29Y82;
  wire tie_high_T29Y82;
  wire tie_low_T30Y82;
  wire tie_high_T30Y82;
  wire tie_low_T31Y82;
  wire tie_high_T31Y82;
  wire tie_low_T32Y82;
  wire tie_high_T32Y82;
  wire tie_low_T33Y82;
  wire tie_high_T33Y82;
  wire tie_low_T34Y82;
  wire tie_high_T34Y82;
  wire tie_low_T35Y82;
  wire tie_high_T35Y82;
  wire tie_low_T0Y83;
  wire tie_high_T0Y83;
  wire tie_low_T1Y83;
  wire tie_high_T1Y83;
  wire tie_low_T2Y83;
  wire tie_high_T2Y83;
  wire tie_low_T3Y83;
  wire tie_high_T3Y83;
  wire tie_low_T4Y83;
  wire tie_high_T4Y83;
  wire tie_low_T5Y83;
  wire tie_high_T5Y83;
  wire tie_low_T6Y83;
  wire tie_high_T6Y83;
  wire tie_low_T7Y83;
  wire tie_high_T7Y83;
  wire tie_low_T8Y83;
  wire tie_high_T8Y83;
  wire tie_low_T9Y83;
  wire tie_high_T9Y83;
  wire tie_low_T10Y83;
  wire tie_high_T10Y83;
  wire tie_low_T11Y83;
  wire tie_high_T11Y83;
  wire tie_low_T12Y83;
  wire tie_high_T12Y83;
  wire tie_low_T13Y83;
  wire tie_high_T13Y83;
  wire tie_low_T14Y83;
  wire tie_high_T14Y83;
  wire tie_low_T15Y83;
  wire tie_high_T15Y83;
  wire tie_low_T16Y83;
  wire tie_high_T16Y83;
  wire tie_low_T17Y83;
  wire tie_high_T17Y83;
  wire tie_low_T18Y83;
  wire tie_high_T18Y83;
  wire tie_low_T19Y83;
  wire tie_high_T19Y83;
  wire tie_low_T20Y83;
  wire tie_high_T20Y83;
  wire tie_low_T21Y83;
  wire tie_high_T21Y83;
  wire tie_low_T22Y83;
  wire tie_high_T22Y83;
  wire tie_low_T23Y83;
  wire tie_high_T23Y83;
  wire tie_low_T24Y83;
  wire tie_high_T24Y83;
  wire tie_low_T25Y83;
  wire tie_high_T25Y83;
  wire tie_low_T26Y83;
  wire tie_high_T26Y83;
  wire tie_low_T27Y83;
  wire tie_high_T27Y83;
  wire tie_low_T28Y83;
  wire tie_high_T28Y83;
  wire tie_low_T29Y83;
  wire tie_high_T29Y83;
  wire tie_low_T30Y83;
  wire tie_high_T30Y83;
  wire tie_low_T31Y83;
  wire tie_high_T31Y83;
  wire tie_low_T32Y83;
  wire tie_high_T32Y83;
  wire tie_low_T33Y83;
  wire tie_high_T33Y83;
  wire tie_low_T34Y83;
  wire tie_high_T34Y83;
  wire tie_low_T35Y83;
  wire tie_high_T35Y83;
  wire tie_low_T0Y84;
  wire tie_high_T0Y84;
  wire tie_low_T1Y84;
  wire tie_high_T1Y84;
  wire tie_low_T2Y84;
  wire tie_high_T2Y84;
  wire tie_low_T3Y84;
  wire tie_high_T3Y84;
  wire tie_low_T4Y84;
  wire tie_high_T4Y84;
  wire tie_low_T5Y84;
  wire tie_high_T5Y84;
  wire tie_low_T6Y84;
  wire tie_high_T6Y84;
  wire tie_low_T7Y84;
  wire tie_high_T7Y84;
  wire tie_low_T8Y84;
  wire tie_high_T8Y84;
  wire tie_low_T9Y84;
  wire tie_high_T9Y84;
  wire tie_low_T10Y84;
  wire tie_high_T10Y84;
  wire tie_low_T11Y84;
  wire tie_high_T11Y84;
  wire tie_low_T12Y84;
  wire tie_high_T12Y84;
  wire tie_low_T13Y84;
  wire tie_high_T13Y84;
  wire tie_low_T14Y84;
  wire tie_high_T14Y84;
  wire tie_low_T15Y84;
  wire tie_high_T15Y84;
  wire tie_low_T16Y84;
  wire tie_high_T16Y84;
  wire tie_low_T17Y84;
  wire tie_high_T17Y84;
  wire tie_low_T18Y84;
  wire tie_high_T18Y84;
  wire tie_low_T19Y84;
  wire tie_high_T19Y84;
  wire tie_low_T20Y84;
  wire tie_high_T20Y84;
  wire tie_low_T21Y84;
  wire tie_high_T21Y84;
  wire tie_low_T22Y84;
  wire tie_high_T22Y84;
  wire tie_low_T23Y84;
  wire tie_high_T23Y84;
  wire tie_low_T24Y84;
  wire tie_high_T24Y84;
  wire tie_low_T25Y84;
  wire tie_high_T25Y84;
  wire tie_low_T26Y84;
  wire tie_high_T26Y84;
  wire tie_low_T27Y84;
  wire tie_high_T27Y84;
  wire tie_low_T28Y84;
  wire tie_high_T28Y84;
  wire tie_low_T29Y84;
  wire tie_high_T29Y84;
  wire tie_low_T30Y84;
  wire tie_high_T30Y84;
  wire tie_low_T31Y84;
  wire tie_high_T31Y84;
  wire tie_low_T32Y84;
  wire tie_high_T32Y84;
  wire tie_low_T33Y84;
  wire tie_high_T33Y84;
  wire tie_low_T34Y84;
  wire tie_high_T34Y84;
  wire tie_low_T35Y84;
  wire tie_high_T35Y84;
  wire tie_low_T0Y85;
  wire tie_high_T0Y85;
  wire tie_low_T1Y85;
  wire tie_high_T1Y85;
  wire tie_low_T2Y85;
  wire tie_high_T2Y85;
  wire tie_low_T3Y85;
  wire tie_high_T3Y85;
  wire tie_low_T4Y85;
  wire tie_high_T4Y85;
  wire tie_low_T5Y85;
  wire tie_high_T5Y85;
  wire tie_low_T6Y85;
  wire tie_high_T6Y85;
  wire tie_low_T7Y85;
  wire tie_high_T7Y85;
  wire tie_low_T8Y85;
  wire tie_high_T8Y85;
  wire tie_low_T9Y85;
  wire tie_high_T9Y85;
  wire tie_low_T10Y85;
  wire tie_high_T10Y85;
  wire tie_low_T11Y85;
  wire tie_high_T11Y85;
  wire tie_low_T12Y85;
  wire tie_high_T12Y85;
  wire tie_low_T13Y85;
  wire tie_high_T13Y85;
  wire tie_low_T14Y85;
  wire tie_high_T14Y85;
  wire tie_low_T15Y85;
  wire tie_high_T15Y85;
  wire tie_low_T16Y85;
  wire tie_high_T16Y85;
  wire tie_low_T17Y85;
  wire tie_high_T17Y85;
  wire tie_low_T18Y85;
  wire tie_high_T18Y85;
  wire tie_low_T19Y85;
  wire tie_high_T19Y85;
  wire tie_low_T20Y85;
  wire tie_high_T20Y85;
  wire tie_low_T21Y85;
  wire tie_high_T21Y85;
  wire tie_low_T22Y85;
  wire tie_high_T22Y85;
  wire tie_low_T23Y85;
  wire tie_high_T23Y85;
  wire tie_low_T24Y85;
  wire tie_high_T24Y85;
  wire tie_low_T25Y85;
  wire tie_high_T25Y85;
  wire tie_low_T26Y85;
  wire tie_high_T26Y85;
  wire tie_low_T27Y85;
  wire tie_high_T27Y85;
  wire tie_low_T28Y85;
  wire tie_high_T28Y85;
  wire tie_low_T29Y85;
  wire tie_high_T29Y85;
  wire tie_low_T30Y85;
  wire tie_high_T30Y85;
  wire tie_low_T31Y85;
  wire tie_high_T31Y85;
  wire tie_low_T32Y85;
  wire tie_high_T32Y85;
  wire tie_low_T33Y85;
  wire tie_high_T33Y85;
  wire tie_low_T34Y85;
  wire tie_high_T34Y85;
  wire tie_low_T35Y85;
  wire tie_high_T35Y85;
  wire tie_low_T0Y86;
  wire tie_high_T0Y86;
  wire tie_low_T1Y86;
  wire tie_high_T1Y86;
  wire tie_low_T2Y86;
  wire tie_high_T2Y86;
  wire tie_low_T3Y86;
  wire tie_high_T3Y86;
  wire tie_low_T4Y86;
  wire tie_high_T4Y86;
  wire tie_low_T5Y86;
  wire tie_high_T5Y86;
  wire tie_low_T6Y86;
  wire tie_high_T6Y86;
  wire tie_low_T7Y86;
  wire tie_high_T7Y86;
  wire tie_low_T8Y86;
  wire tie_high_T8Y86;
  wire tie_low_T9Y86;
  wire tie_high_T9Y86;
  wire tie_low_T10Y86;
  wire tie_high_T10Y86;
  wire tie_low_T11Y86;
  wire tie_high_T11Y86;
  wire tie_low_T12Y86;
  wire tie_high_T12Y86;
  wire tie_low_T13Y86;
  wire tie_high_T13Y86;
  wire tie_low_T14Y86;
  wire tie_high_T14Y86;
  wire tie_low_T15Y86;
  wire tie_high_T15Y86;
  wire tie_low_T16Y86;
  wire tie_high_T16Y86;
  wire tie_low_T17Y86;
  wire tie_high_T17Y86;
  wire tie_low_T18Y86;
  wire tie_high_T18Y86;
  wire tie_low_T19Y86;
  wire tie_high_T19Y86;
  wire tie_low_T20Y86;
  wire tie_high_T20Y86;
  wire tie_low_T21Y86;
  wire tie_high_T21Y86;
  wire tie_low_T22Y86;
  wire tie_high_T22Y86;
  wire tie_low_T23Y86;
  wire tie_high_T23Y86;
  wire tie_low_T24Y86;
  wire tie_high_T24Y86;
  wire tie_low_T25Y86;
  wire tie_high_T25Y86;
  wire tie_low_T26Y86;
  wire tie_high_T26Y86;
  wire tie_low_T27Y86;
  wire tie_high_T27Y86;
  wire tie_low_T28Y86;
  wire tie_high_T28Y86;
  wire tie_low_T29Y86;
  wire tie_high_T29Y86;
  wire tie_low_T30Y86;
  wire tie_high_T30Y86;
  wire tie_low_T31Y86;
  wire tie_high_T31Y86;
  wire tie_low_T32Y86;
  wire tie_high_T32Y86;
  wire tie_low_T33Y86;
  wire tie_high_T33Y86;
  wire tie_low_T34Y86;
  wire tie_high_T34Y86;
  wire tie_low_T35Y86;
  wire tie_high_T35Y86;
  wire tie_low_T0Y87;
  wire tie_high_T0Y87;
  wire tie_low_T1Y87;
  wire tie_high_T1Y87;
  wire tie_low_T2Y87;
  wire tie_high_T2Y87;
  wire tie_low_T3Y87;
  wire tie_high_T3Y87;
  wire tie_low_T4Y87;
  wire tie_high_T4Y87;
  wire tie_low_T5Y87;
  wire tie_high_T5Y87;
  wire tie_low_T6Y87;
  wire tie_high_T6Y87;
  wire tie_low_T7Y87;
  wire tie_high_T7Y87;
  wire tie_low_T8Y87;
  wire tie_high_T8Y87;
  wire tie_low_T9Y87;
  wire tie_high_T9Y87;
  wire tie_low_T10Y87;
  wire tie_high_T10Y87;
  wire tie_low_T11Y87;
  wire tie_high_T11Y87;
  wire tie_low_T12Y87;
  wire tie_high_T12Y87;
  wire tie_low_T13Y87;
  wire tie_high_T13Y87;
  wire tie_low_T14Y87;
  wire tie_high_T14Y87;
  wire tie_low_T15Y87;
  wire tie_high_T15Y87;
  wire tie_low_T16Y87;
  wire tie_high_T16Y87;
  wire tie_low_T17Y87;
  wire tie_high_T17Y87;
  wire tie_low_T18Y87;
  wire tie_high_T18Y87;
  wire tie_low_T19Y87;
  wire tie_high_T19Y87;
  wire tie_low_T20Y87;
  wire tie_high_T20Y87;
  wire tie_low_T21Y87;
  wire tie_high_T21Y87;
  wire tie_low_T22Y87;
  wire tie_high_T22Y87;
  wire tie_low_T23Y87;
  wire tie_high_T23Y87;
  wire tie_low_T24Y87;
  wire tie_high_T24Y87;
  wire tie_low_T25Y87;
  wire tie_high_T25Y87;
  wire tie_low_T26Y87;
  wire tie_high_T26Y87;
  wire tie_low_T27Y87;
  wire tie_high_T27Y87;
  wire tie_low_T28Y87;
  wire tie_high_T28Y87;
  wire tie_low_T29Y87;
  wire tie_high_T29Y87;
  wire tie_low_T30Y87;
  wire tie_high_T30Y87;
  wire tie_low_T31Y87;
  wire tie_high_T31Y87;
  wire tie_low_T32Y87;
  wire tie_high_T32Y87;
  wire tie_low_T33Y87;
  wire tie_high_T33Y87;
  wire tie_low_T34Y87;
  wire tie_high_T34Y87;
  wire tie_low_T35Y87;
  wire tie_high_T35Y87;
  wire tie_low_T0Y88;
  wire tie_high_T0Y88;
  wire tie_low_T1Y88;
  wire tie_high_T1Y88;
  wire tie_low_T2Y88;
  wire tie_high_T2Y88;
  wire tie_low_T3Y88;
  wire tie_high_T3Y88;
  wire tie_low_T4Y88;
  wire tie_high_T4Y88;
  wire tie_low_T5Y88;
  wire tie_high_T5Y88;
  wire tie_low_T6Y88;
  wire tie_high_T6Y88;
  wire tie_low_T7Y88;
  wire tie_high_T7Y88;
  wire tie_low_T8Y88;
  wire tie_high_T8Y88;
  wire tie_low_T9Y88;
  wire tie_high_T9Y88;
  wire tie_low_T10Y88;
  wire tie_high_T10Y88;
  wire tie_low_T11Y88;
  wire tie_high_T11Y88;
  wire tie_low_T12Y88;
  wire tie_high_T12Y88;
  wire tie_low_T13Y88;
  wire tie_high_T13Y88;
  wire tie_low_T14Y88;
  wire tie_high_T14Y88;
  wire tie_low_T15Y88;
  wire tie_high_T15Y88;
  wire tie_low_T16Y88;
  wire tie_high_T16Y88;
  wire tie_low_T17Y88;
  wire tie_high_T17Y88;
  wire tie_low_T18Y88;
  wire tie_high_T18Y88;
  wire tie_low_T19Y88;
  wire tie_high_T19Y88;
  wire tie_low_T20Y88;
  wire tie_high_T20Y88;
  wire tie_low_T21Y88;
  wire tie_high_T21Y88;
  wire tie_low_T22Y88;
  wire tie_high_T22Y88;
  wire tie_low_T23Y88;
  wire tie_high_T23Y88;
  wire tie_low_T24Y88;
  wire tie_high_T24Y88;
  wire tie_low_T25Y88;
  wire tie_high_T25Y88;
  wire tie_low_T26Y88;
  wire tie_high_T26Y88;
  wire tie_low_T27Y88;
  wire tie_high_T27Y88;
  wire tie_low_T28Y88;
  wire tie_high_T28Y88;
  wire tie_low_T29Y88;
  wire tie_high_T29Y88;
  wire tie_low_T30Y88;
  wire tie_high_T30Y88;
  wire tie_low_T31Y88;
  wire tie_high_T31Y88;
  wire tie_low_T32Y88;
  wire tie_high_T32Y88;
  wire tie_low_T33Y88;
  wire tie_high_T33Y88;
  wire tie_low_T34Y88;
  wire tie_high_T34Y88;
  wire tie_low_T35Y88;
  wire tie_high_T35Y88;
  wire tie_low_T0Y89;
  wire tie_high_T0Y89;
  wire tie_low_T1Y89;
  wire tie_high_T1Y89;
  wire tie_low_T2Y89;
  wire tie_high_T2Y89;
  wire tie_low_T3Y89;
  wire tie_high_T3Y89;
  wire tie_low_T4Y89;
  wire tie_high_T4Y89;
  wire tie_low_T5Y89;
  wire tie_high_T5Y89;
  wire tie_low_T6Y89;
  wire tie_high_T6Y89;
  wire tie_low_T7Y89;
  wire tie_high_T7Y89;
  wire tie_low_T8Y89;
  wire tie_high_T8Y89;
  wire tie_low_T9Y89;
  wire tie_high_T9Y89;
  wire tie_low_T10Y89;
  wire tie_high_T10Y89;
  wire tie_low_T11Y89;
  wire tie_high_T11Y89;
  wire tie_low_T12Y89;
  wire tie_high_T12Y89;
  wire tie_low_T13Y89;
  wire tie_high_T13Y89;
  wire tie_low_T14Y89;
  wire tie_high_T14Y89;
  wire tie_low_T15Y89;
  wire tie_high_T15Y89;
  wire tie_low_T16Y89;
  wire tie_high_T16Y89;
  wire tie_low_T17Y89;
  wire tie_high_T17Y89;
  wire tie_low_T18Y89;
  wire tie_high_T18Y89;
  wire tie_low_T19Y89;
  wire tie_high_T19Y89;
  wire tie_low_T20Y89;
  wire tie_high_T20Y89;
  wire tie_low_T21Y89;
  wire tie_high_T21Y89;
  wire tie_low_T22Y89;
  wire tie_high_T22Y89;
  wire tie_low_T23Y89;
  wire tie_high_T23Y89;
  wire tie_low_T24Y89;
  wire tie_high_T24Y89;
  wire tie_low_T25Y89;
  wire tie_high_T25Y89;
  wire tie_low_T26Y89;
  wire tie_high_T26Y89;
  wire tie_low_T27Y89;
  wire tie_high_T27Y89;
  wire tie_low_T28Y89;
  wire tie_high_T28Y89;
  wire tie_low_T29Y89;
  wire tie_high_T29Y89;
  wire tie_low_T30Y89;
  wire tie_high_T30Y89;
  wire tie_low_T31Y89;
  wire tie_high_T31Y89;
  wire tie_low_T32Y89;
  wire tie_high_T32Y89;
  wire tie_low_T33Y89;
  wire tie_high_T33Y89;
  wire tie_low_T34Y89;
  wire tie_high_T34Y89;
  wire tie_low_T35Y89;
  wire tie_high_T35Y89;

  // Cell instances
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10000  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(126));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10001  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(128));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10002  (.A(128), .Y(129));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10003  (.A(tie_low_T4Y41), .B(tie_low_T4Y41), .Y(131));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10004  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(133));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10005  (.A(133), .Y(134));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10006  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(135));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10007  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(136));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10008  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(137));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10009  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(139));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10010  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(140));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10011  (.A(140), .Y(141));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10012  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .Y(144));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10013  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(147));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10014  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(149));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10015  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(151));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10016  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(154));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10017  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(155));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10018  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(156));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10019  (.A(156), .Y(157));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10020  (.A(tie_low_T4Y40), .B(tie_low_T4Y40), .Y(158));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10021  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(159));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10022  (.A(159), .Y(160));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10023  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .X(161));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10024  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(162));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10025  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(163));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10026  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(164));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10027  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(165));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10028  (.A(165), .Y(166));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10029  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(168));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10030  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(170));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10031  (.A(tie_low_T6Y17), .B(tie_low_T6Y17), .X(173));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10032  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(174));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10033  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .Y(176));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10034  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(177));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10035  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(178));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10036  (.A(178), .Y(179));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10037  (.A(tie_low_T5Y37), .B(tie_low_T5Y37), .Y(180));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10038  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(181));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10039  (.A(181), .Y(182));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10040  (.A(tie_low_T2Y45), .B(tie_low_T2Y45), .X(183));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10041  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(184));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10042  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(185));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10043  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(186));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10044  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(187));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10045  (.A(187), .Y(188));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10046  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .Y(190));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10047  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(192));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10048  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(193));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10049  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(195));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10050  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(196));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10051  (.A(196), .Y(197));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10052  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(198));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10053  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(200));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10054  (.A(200), .Y(201));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10055  (.A(tie_low_T4Y40), .B(tie_low_T4Y40), .Y(202));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10056  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(203));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10057  (.A(203), .Y(204));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10058  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .X(205));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10059  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(206));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10060  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(207));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10061  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(208));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10062  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(209));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10063  (.A(209), .Y(210));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10064  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(212));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10065  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(214));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10066  (.A(tie_low_T6Y17), .B(tie_low_T6Y17), .X(216));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10067  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(217));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10068  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(219));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10069  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(220));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10070  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(221));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10071  (.A(221), .Y(222));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10072  (.A(tie_low_T4Y40), .B(tie_low_T4Y40), .Y(223));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10073  (.A(tie_low_T1Y47), .B(tie_low_T1Y47), .Y(224));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10074  (.A(224), .Y(225));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10075  (.A(tie_low_T0Y47), .B(tie_low_T0Y47), .X(226));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10076  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(227));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10077  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(228));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10078  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(229));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10079  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(230));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10080  (.A(230), .Y(231));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10081  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .Y(233));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10082  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .Y(235));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10083  (.A(tie_low_T6Y17), .B(tie_low_T6Y17), .X(237));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10084  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(238));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10085  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(240));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10086  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(241));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10087  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(242));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10088  (.A(242), .Y(243));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10089  (.A(tie_low_T4Y39), .B(tie_low_T4Y39), .Y(244));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10090  (.A(tie_low_T1Y46), .B(tie_low_T1Y46), .Y(245));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10091  (.A(245), .Y(246));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10092  (.A(tie_low_T1Y47), .B(tie_low_T1Y47), .X(247));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10093  (.A(tie_low_T1Y47), .B(tie_low_T1Y47), .Y(248));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10094  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(249));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10095  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(250));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10096  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(251));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10097  (.A(251), .Y(252));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10098  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(255));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10099  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(257));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10100  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(259));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10101  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(260));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10102  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(261));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10103  (.A(261), .Y(262));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10104  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(265));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10105  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(266));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10106  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .Y(267));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10107  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(268));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10108  (.A(268), .Y(269));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10109  (.A(tie_low_T6Y35), .B(tie_low_T6Y35), .Y(270));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10110  (.A(tie_low_T1Y46), .B(tie_low_T1Y46), .Y(271));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10111  (.A(271), .Y(272));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10112  (.A(tie_low_T3Y43), .B(tie_low_T3Y43), .X(273));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10113  (.A(tie_low_T1Y47), .B(tie_low_T1Y47), .Y(274));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10114  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(275));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10115  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(276));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10116  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(277));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10117  (.A(277), .Y(278));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10118  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(280));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10119  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(282));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10120  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(284));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10121  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(285));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10122  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(288));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10123  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(289));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10124  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(290));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10125  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(291));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10126  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(292));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10127  (.A(292), .Y(293));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10128  (.A(tie_low_T6Y35), .B(tie_low_T6Y35), .Y(294));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10129  (.A(tie_low_T1Y46), .B(tie_low_T1Y46), .Y(295));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10130  (.A(295), .Y(296));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10131  (.A(tie_low_T3Y43), .B(tie_low_T3Y43), .X(297));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10132  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(298));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10133  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(299));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10134  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(300));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10135  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(301));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10136  (.A(301), .Y(302));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10137  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(304));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10138  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .Y(306));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10139  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .Y(308));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10140  (.A(tie_low_T8Y21), .B(tie_low_T8Y21), .X(310));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10141  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(311));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10142  (.A(311), .Y(312));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10143  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(313));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10144  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(314));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10145  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(315));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10146  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(316));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10147  (.A(316), .Y(317));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10148  (.A(tie_low_T6Y36), .B(tie_low_T6Y36), .Y(318));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10149  (.A(tie_low_T1Y47), .B(tie_low_T1Y47), .Y(319));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10150  (.A(319), .Y(320));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10151  (.A(tie_low_T2Y44), .B(tie_low_T2Y44), .X(321));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10152  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(322));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10153  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(323));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10154  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(324));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10155  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(325));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10156  (.A(325), .Y(326));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10157  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(328));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10158  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(330));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10159  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(332));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10160  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(333));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10161  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(334));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10162  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(335));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10163  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(336));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10164  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(337));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10165  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(338));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10166  (.A(338), .Y(339));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10167  (.A(tie_low_T6Y36), .B(tie_low_T6Y36), .Y(340));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10168  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(341));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10169  (.A(341), .Y(342));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10170  (.A(tie_low_T2Y44), .B(tie_low_T2Y44), .X(343));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10171  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(344));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10172  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(345));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10173  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(346));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10174  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(347));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10175  (.A(347), .Y(348));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10176  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(350));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10177  (.A(350), .Y(351));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10178  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(353));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10179  (.A(353), .Y(354));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10180  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(356));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10181  (.A(tie_low_T8Y20), .B(tie_low_T8Y20), .X(357));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10182  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(358));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10183  (.A(358), .Y(359));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10184  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(360));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10185  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(361));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10186  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(362));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10187  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(363));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10188  (.A(tie_low_T5Y34), .B(tie_low_T5Y34), .X(364));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10189  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(365));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10190  (.A(365), .Y(366));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10191  (.A(tie_low_T2Y45), .B(tie_low_T2Y45), .X(367));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10192  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(368));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10193  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(369));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10194  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(370));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10195  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(371));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10196  (.A(371), .Y(372));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10197  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(374));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10198  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(376));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10199  (.A(376), .Y(377));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10200  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(379));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10201  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(380));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10202  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(381));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10203  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(382));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10204  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(383));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10205  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(384));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10206  (.A(384), .Y(385));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10207  (.A(tie_low_T6Y37), .B(tie_low_T6Y37), .Y(386));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10208  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(387));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10209  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(388));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10210  (.A(388), .Y(389));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10211  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .X(390));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10212  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(391));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10213  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(392));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10214  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(393));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10215  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(394));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10216  (.A(394), .Y(395));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10217  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(397));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10218  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(399));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10219  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(401));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10220  (.A(tie_low_T8Y20), .B(tie_low_T8Y20), .X(402));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10221  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(403));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10222  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(404));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10223  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(405));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10224  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(406));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10225  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(407));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10226  (.A(407), .Y(408));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10227  (.A(tie_low_T5Y38), .B(tie_low_T5Y38), .Y(409));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10228  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(410));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10229  (.A(tie_low_T1Y47), .B(tie_low_T1Y47), .X(411));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10230  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(412));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10231  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(413));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10232  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(414));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10233  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(415));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10234  (.A(415), .Y(416));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10235  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(418));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10236  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(420));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10237  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(422));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10238  (.A(tie_low_T8Y21), .B(tie_low_T8Y21), .X(423));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10239  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(424));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10240  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(425));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10241  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(426));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10242  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(427));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10243  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(428));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10244  (.A(428), .Y(429));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10245  (.A(tie_low_T5Y44), .B(tie_low_T5Y44), .Y(430));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10246  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(431));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10247  (.A(tie_low_T0Y52), .B(tie_low_T0Y52), .Y(432));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10248  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(434));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10249  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(435));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10250  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(436));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10251  (.A(tie_low_T13Y39), .B(tie_low_T13Y39), .Y(437));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10252  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(439));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10253  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(441));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10254  (.A(tie_low_T13Y39), .B(tie_low_T13Y39), .Y(442));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10255  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(444));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10256  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(446));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10257  (.A(tie_low_T13Y39), .B(tie_low_T13Y39), .Y(447));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10258  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(449));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10259  (.A(tie_low_T0Y50), .B(tie_low_T0Y50), .Y(451));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10260  (.A(tie_low_T13Y39), .B(tie_low_T13Y39), .Y(452));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10261  (.A(tie_low_T21Y24), .B(tie_low_T21Y24), .X(455));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10262  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(457));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10263  (.A(tie_low_T35Y60), .B(tie_low_T35Y60), .Y(458));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10264  (.A(tie_low_T21Y31), .B(tie_low_T21Y31), .Y(460));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10265  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(461));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10266  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(463));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10267  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(464));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10268  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(465));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10269  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(467));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10270  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(470));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10271  (.A(470), .Y(471));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10272  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .Y(473));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10273  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(475));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10274  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(477));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10275  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(478));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10276  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(479));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10277  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .X(480));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10278  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(483));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10279  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(485));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10280  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(486));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10281  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(487));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10282  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .X(490));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10283  (.A(490), .Y(491));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10284  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(492));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10285  (.A(492), .Y(493));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10286  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(495));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10287  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .X(497));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10288  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(498));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10289  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .X(499));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10290  (.A(tie_low_T13Y22), .B(tie_low_T13Y22), .Y(500));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10291  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(502));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10292  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(503));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10293  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .Y(504));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10294  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(505));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10295  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(506));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10296  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(507));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10297  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(509));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10298  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(510));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10299  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .X(512));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10300  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(513));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10301  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(514));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10302  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(515));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10303  (.A(tie_low_T8Y25), .B(tie_low_T8Y25), .X(517));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10304  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(519));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10305  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(520));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10306  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(521));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10307  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(522));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10308  (.A(522), .Y(523));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10309  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(524));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10310  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(525));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10311  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(526));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10312  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(527));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10313  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(528));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10314  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(529));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10315  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(530));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10316  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .Y(532));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10317  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(533));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10318  (.A(533), .Y(534));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10319  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(535));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10320  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(536));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10321  (.A(536), .Y(537));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10322  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(538));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10323  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(540));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10324  (.A(540), .Y(541));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10325  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .Y(543));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10326  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .X(545));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10327  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .X(547));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10328  (.A(547), .Y(548));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10329  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .Y(549));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10330  (.A(tie_low_T12Y27), .B(tie_low_T12Y27), .X(551));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10331  (.A(tie_low_T35Y60), .B(tie_low_T35Y60), .Y(553));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10332  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(555));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10333  (.A(tie_low_T15Y18), .B(tie_low_T15Y18), .X(556));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10334  (.A(tie_low_T9Y12), .B(tie_low_T9Y12), .Y(557));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10335  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(558));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10336  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(559));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10337  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .Y(560));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10338  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(561));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10339  (.A(tie_low_T11Y15), .B(tie_low_T11Y15), .Y(563));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10340  (.A(563), .Y(564));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10341  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(565));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10342  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(566));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10343  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(568));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10344  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .Y(569));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10345  (.A(569), .Y(570));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10346  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .Y(571));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10347  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(572));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10348  (.A(tie_low_T11Y11), .B(tie_low_T11Y11), .X(573));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10349  (.A(tie_low_T20Y26), .B(tie_low_T20Y26), .X(574));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10350  (.A(tie_low_T16Y17), .B(tie_low_T16Y17), .X(575));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10351  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(576));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10352  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(578));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10353  (.A(578), .Y(579));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10354  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(580));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10355  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .X(581));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10356  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(582));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10357  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(584));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10358  (.A(tie_low_T16Y50), .B(tie_low_T16Y50), .Y(586));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10359  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .X(589));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10360  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(591));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10361  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(592));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10362  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(594));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10363  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .X(596));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10364  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(598));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10365  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(599));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10366  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(601));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10367  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(602));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10368  (.A(tie_low_T9Y14), .B(tie_low_T9Y14), .Y(604));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10369  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(607));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10370  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(610));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10371  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(612));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10372  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(613));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10373  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(616));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10374  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(618));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10375  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(619));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10376  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(620));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10377  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(622));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10378  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(624));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10379  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(625));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10380  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(626));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10381  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(627));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10382  (.A(627), .Y(628));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10383  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .Y(630));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10384  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(632));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10385  (.A(632), .Y(633));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10386  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(635));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10387  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(636));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10388  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .X(637));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10389  (.A(637), .Y(638));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10390  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(640));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10391  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(643));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10392  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(644));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10393  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(645));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10394  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(646));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10395  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(647));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10396  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(648));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10397  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .X(649));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10398  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .X(651));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10399  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .X(652));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10400  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(653));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10401  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(655));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10402  (.A(655), .Y(656));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10403  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(657));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10404  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .Y(658));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10405  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(659));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10406  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(660));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10407  (.A(660), .Y(661));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10408  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(662));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10409  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .Y(663));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10410  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(664));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10411  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(665));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10412  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(667));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10413  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(668));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10414  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .Y(669));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10415  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .X(670));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10416  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .X(671));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10417  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(672));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10418  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .X(673));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10419  (.A(673), .Y(674));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10420  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .Y(676));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10421  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(677));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10422  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(679));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10423  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(680));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10424  (.A(tie_low_T10Y16), .B(tie_low_T10Y16), .Y(682));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10425  (.A(682), .Y(683));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10426  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(684));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10427  (.A(684), .Y(685));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10428  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(686));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10429  (.A(686), .Y(687));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10430  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .Y(688));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10431  (.A(688), .Y(689));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10432  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(84));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10433  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .Y(692));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10434  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(693));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10435  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(695));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10436  (.A(695), .Y(696));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10437  (.A(tie_low_T10Y32), .B(tie_low_T10Y32), .X(698));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10438  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(699));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10439  (.A(tie_low_T16Y13), .B(tie_low_T16Y13), .X(700));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10440  (.A(700), .Y(701));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10441  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(702));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10442  (.A(tie_low_T17Y11), .B(tie_low_T17Y11), .Y(703));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10443  (.A(tie_low_T11Y3), .B(tie_low_T11Y3), .Y(704));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10444  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(706));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10445  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .X(708));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10446  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(709));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10447  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(710));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10448  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(712));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10449  (.A(712), .Y(713));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10450  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(716));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10451  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(717));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10452  (.A(tie_low_T11Y30), .B(tie_low_T11Y30), .X(718));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10453  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(720));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10454  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(722));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10455  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(723));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10456  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(725));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10457  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(726));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10458  (.A(tie_low_T14Y14), .B(tie_low_T14Y14), .Y(727));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10459  (.A(tie_low_T12Y25), .B(tie_low_T12Y25), .Y(728));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10460  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .X(730));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10461  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .X(731));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10462  (.A(731), .Y(732));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10463  (.A(tie_low_T3Y0), .B(tie_low_T3Y0), .Y(85));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10464  (.A(tie_low_T3Y0), .B(tie_low_T3Y0), .Y(733));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10465  (.A(tie_low_T17Y10), .B(tie_low_T17Y10), .Y(734));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10466  (.A(tie_low_T13Y3), .B(tie_low_T13Y3), .Y(735));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10467  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(738));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10468  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(740));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10469  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(741));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10470  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(742));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10471  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(744));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10472  (.A(744), .Y(745));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10473  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(747));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10474  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(748));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10475  (.A(tie_low_T11Y31), .B(tie_low_T11Y31), .X(749));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10476  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(750));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10477  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .Y(751));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10478  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(752));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10479  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(754));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10480  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(755));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10481  (.A(tie_low_T14Y14), .B(tie_low_T14Y14), .Y(756));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10482  (.A(tie_low_T14Y14), .B(tie_low_T14Y14), .X(757));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10483  (.A(757), .Y(758));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10484  (.A(tie_low_T9Y27), .B(tie_low_T9Y27), .Y(759));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10485  (.A(759), .Y(760));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10486  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .Y(761));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10487  (.A(761), .Y(762));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10488  (.A(tie_low_T7Y0), .B(tie_low_T7Y0), .Y(86));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10489  (.A(tie_low_T7Y0), .B(tie_low_T7Y0), .Y(763));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10490  (.A(tie_low_T17Y11), .B(tie_low_T17Y11), .Y(764));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10491  (.A(tie_low_T14Y3), .B(tie_low_T14Y3), .Y(765));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10492  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(767));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10493  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(769));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10494  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(770));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10495  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(771));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10496  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(773));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10497  (.A(773), .Y(774));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10498  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(776));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10499  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(777));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10500  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .X(778));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10501  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(779));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10502  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(780));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10503  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(781));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10504  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(782));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10505  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(783));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10506  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(784));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10507  (.A(784), .Y(785));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10508  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(786));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10509  (.A(786), .Y(787));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10510  (.A(tie_low_T9Y27), .B(tie_low_T9Y27), .Y(788));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10511  (.A(788), .Y(789));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10512  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(790));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10513  (.A(790), .Y(791));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10514  (.A(tie_low_T11Y0), .B(tie_low_T11Y0), .Y(87));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10515  (.A(tie_low_T17Y11), .B(tie_low_T17Y11), .Y(792));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10516  (.A(tie_low_T11Y0), .B(tie_low_T11Y0), .Y(793));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10517  (.A(tie_low_T15Y3), .B(tie_low_T15Y3), .Y(794));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10518  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(796));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10519  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(798));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10520  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(799));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10521  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(800));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10522  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .X(802));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10523  (.A(802), .Y(803));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10524  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(805));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10525  (.A(tie_low_T13Y20), .B(tie_low_T13Y20), .Y(806));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10526  (.A(tie_low_T13Y31), .B(tie_low_T13Y31), .X(807));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10527  (.A(tie_low_T13Y20), .B(tie_low_T13Y20), .X(808));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10528  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(809));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10529  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(810));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10530  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(811));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10531  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(812));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10532  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(813));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10533  (.A(813), .Y(814));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10534  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .Y(815));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10535  (.A(815), .Y(816));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10536  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(817));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10537  (.A(817), .Y(818));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10538  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(819));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10539  (.A(819), .Y(820));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10540  (.A(tie_low_T15Y0), .B(tie_low_T15Y0), .Y(88));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10541  (.A(tie_low_T15Y0), .B(tie_low_T15Y0), .Y(821));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10542  (.A(tie_low_T17Y10), .B(tie_low_T17Y10), .Y(822));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10543  (.A(tie_low_T17Y3), .B(tie_low_T17Y3), .Y(823));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10544  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(825));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10545  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(827));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10546  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(828));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10547  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .X(829));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10548  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .X(831));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10549  (.A(831), .Y(832));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10550  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(834));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10551  (.A(tie_low_T13Y20), .B(tie_low_T13Y20), .Y(835));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10552  (.A(tie_low_T13Y31), .B(tie_low_T13Y31), .X(836));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10553  (.A(tie_low_T13Y20), .B(tie_low_T13Y20), .X(837));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10554  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .Y(838));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10555  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(839));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10556  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(840));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10557  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(841));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10558  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(842));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10559  (.A(842), .Y(843));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10560  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(844));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10561  (.A(844), .Y(845));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10562  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(846));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10563  (.A(846), .Y(847));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10564  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .Y(848));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10565  (.A(848), .Y(849));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10566  (.A(tie_low_T19Y0), .B(tie_low_T19Y0), .Y(89));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10567  (.A(tie_low_T19Y0), .B(tie_low_T19Y0), .Y(850));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10568  (.A(tie_low_T17Y11), .B(tie_low_T17Y11), .Y(851));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10569  (.A(tie_low_T18Y4), .B(tie_low_T18Y4), .Y(852));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10570  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(854));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10571  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(856));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10572  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(857));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10573  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(858));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10574  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(860));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10575  (.A(860), .Y(861));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10576  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(863));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10577  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(864));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10578  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .X(865));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10579  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .X(866));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10580  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(867));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10581  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(868));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10582  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(869));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10583  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(870));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10584  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(871));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10585  (.A(871), .Y(872));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10586  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(873));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10587  (.A(873), .Y(874));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10588  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(875));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10589  (.A(875), .Y(876));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10590  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(877));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10591  (.A(877), .Y(878));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10592  (.A(tie_low_T23Y0), .B(tie_low_T23Y0), .Y(90));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10593  (.A(tie_low_T17Y11), .B(tie_low_T17Y11), .Y(879));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10594  (.A(tie_low_T23Y0), .B(tie_low_T23Y0), .Y(880));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10595  (.A(tie_low_T19Y4), .B(tie_low_T19Y4), .Y(881));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10596  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(883));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10597  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(885));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10598  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(886));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10599  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .X(887));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10600  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .X(889));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10601  (.A(889), .Y(890));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10602  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(892));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10603  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(893));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10604  (.A(tie_low_T9Y27), .B(tie_low_T9Y27), .X(894));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10605  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .X(895));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10606  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(896));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10607  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .Y(897));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10608  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(898));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10609  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .Y(899));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10610  (.A(899), .Y(900));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10611  (.A(tie_low_T14Y14), .B(tie_low_T14Y14), .Y(901));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10612  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(902));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10613  (.A(902), .Y(903));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10614  (.A(tie_low_T16Y25), .B(tie_low_T16Y25), .Y(904));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10615  (.A(tie_low_T22Y12), .B(tie_low_T22Y12), .X(905));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10616  (.A(tie_low_T27Y0), .B(tie_low_T27Y0), .X(91));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10617  (.A(tie_low_T27Y0), .B(tie_low_T27Y0), .Y(906));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10618  (.A(tie_low_T17Y11), .B(tie_low_T17Y11), .Y(907));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10619  (.A(tie_low_T21Y4), .B(tie_low_T21Y4), .Y(908));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10620  (.A(tie_low_T17Y22), .B(tie_low_T17Y22), .Y(909));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10621  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(910));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10622  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(911));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10623  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(912));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10624  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(913));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10625  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(914));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10626  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(915));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10627  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(916));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10628  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(917));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10629  (.A(917), .Y(918));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10630  (.A(tie_low_T31Y0), .B(tie_low_T31Y0), .Y(92));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10631  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(919));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10632  (.A(tie_low_T31Y0), .B(tie_low_T31Y0), .Y(920));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10633  (.A(tie_low_T22Y4), .B(tie_low_T22Y4), .Y(921));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10634  (.A(tie_low_T17Y20), .B(tie_low_T17Y20), .Y(922));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10635  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(923));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10636  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(924));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10637  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(925));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10638  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(926));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10639  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(927));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10640  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .X(928));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10641  (.A(928), .Y(929));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10642  (.A(tie_low_T35Y0), .B(tie_low_T35Y0), .Y(93));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10643  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(930));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10644  (.A(tie_low_T35Y0), .B(tie_low_T35Y0), .Y(931));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10645  (.A(tie_low_T23Y4), .B(tie_low_T23Y4), .Y(932));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10646  (.A(tie_low_T18Y22), .B(tie_low_T18Y22), .Y(933));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10647  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(934));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10648  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(935));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10649  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(936));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10650  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(937));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10651  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .Y(938));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10652  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(939));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10653  (.A(939), .Y(940));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10654  (.A(tie_low_T35Y0), .B(tie_low_T35Y0), .Y(94));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10655  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(941));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10656  (.A(tie_low_T35Y0), .B(tie_low_T35Y0), .Y(942));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10657  (.A(tie_low_T23Y4), .B(tie_low_T23Y4), .Y(943));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10658  (.A(tie_low_T17Y22), .B(tie_low_T17Y22), .Y(944));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10659  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(945));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10660  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(946));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10661  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(947));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10662  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(948));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10663  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(949));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10664  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(950));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10665  (.A(950), .Y(951));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10666  (.A(tie_low_T35Y10), .B(tie_low_T35Y10), .Y(95));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10667  (.A(tie_low_T35Y10), .B(tie_low_T35Y10), .Y(952));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10668  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(953));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10669  (.A(tie_low_T23Y8), .B(tie_low_T23Y8), .Y(954));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10670  (.A(tie_low_T18Y24), .B(tie_low_T18Y24), .Y(955));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10671  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .Y(956));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10672  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(957));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10673  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(958));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10674  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .Y(959));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10675  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(960));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10676  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(961));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10677  (.A(961), .Y(962));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10678  (.A(tie_low_T35Y20), .B(tie_low_T35Y20), .Y(96));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10679  (.A(tie_low_T35Y20), .B(tie_low_T35Y20), .Y(963));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10680  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(964));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10681  (.A(tie_low_T23Y11), .B(tie_low_T23Y11), .Y(965));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10682  (.A(tie_low_T18Y25), .B(tie_low_T18Y25), .Y(966));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10683  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(967));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10684  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(968));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10685  (.A(tie_low_T9Y26), .B(tie_low_T9Y26), .Y(969));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10686  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(970));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10687  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(971));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10688  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(972));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10689  (.A(972), .Y(973));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10690  (.A(tie_low_T35Y30), .B(tie_low_T35Y30), .Y(97));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10691  (.A(tie_low_T35Y30), .B(tie_low_T35Y30), .Y(974));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10692  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(975));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10693  (.A(tie_low_T23Y14), .B(tie_low_T23Y14), .Y(976));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10694  (.A(tie_low_T17Y30), .B(tie_low_T17Y30), .Y(977));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10695  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(978));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10696  (.A(978), .Y(979));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10697  (.A(213), .B(659), .Y(980));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10698  (.A(980), .Y(981));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10699  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(982));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10700  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(983));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10701  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(984));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10702  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(985));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10703  (.A(985), .Y(986));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10704  (.A(tie_low_T35Y40), .B(tie_low_T35Y40), .Y(98));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10705  (.A(tie_low_T35Y40), .B(tie_low_T35Y40), .Y(987));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10706  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(988));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10707  (.A(tie_low_T23Y18), .B(tie_low_T23Y18), .Y(989));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10708  (.A(tie_low_T21Y31), .B(tie_low_T21Y31), .Y(990));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10709  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .Y(991));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10710  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .Y(992));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10711  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(993));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10712  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .Y(994));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10713  (.A(tie_low_T12Y24), .B(tie_low_T12Y24), .Y(995));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10714  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .X(996));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10715  (.A(996), .Y(997));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10716  (.A(tie_low_T35Y50), .B(tie_low_T35Y50), .Y(99));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10717  (.A(tie_low_T35Y50), .B(tie_low_T35Y50), .Y(998));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10718  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(999));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10719  (.A(tie_low_T23Y21), .B(tie_low_T23Y21), .Y(1000));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10720  (.A(39), .B(695), .Y(1001));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10721  (.A(tie_low_T12Y25), .B(tie_low_T12Y25), .X(1003));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10722  (.A(1003), .Y(1004));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10723  (.A(tie_low_T13Y22), .B(tie_low_T13Y22), .X(1005));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10724  (.A(tie_low_T14Y21), .B(tie_low_T14Y21), .Y(1007));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10725  (.A(tie_low_T15Y15), .B(tie_low_T15Y15), .Y(1008));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10726  (.A(tie_low_T13Y23), .B(tie_low_T13Y23), .X(1009));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10727  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(1011));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10728  (.A(tie_low_T15Y15), .B(tie_low_T15Y15), .Y(1012));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10729  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(1014));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10730  (.A(tie_low_T13Y23), .B(tie_low_T13Y23), .X(1016));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10731  (.A(tie_low_T15Y15), .B(tie_low_T15Y15), .Y(1017));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10732  (.A(tie_low_T13Y24), .B(tie_low_T13Y24), .X(1018));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10733  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(1020));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10734  (.A(tie_low_T15Y15), .B(tie_low_T15Y15), .Y(1021));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10735  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .Y(1022));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10736  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(1024));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10737  (.A(tie_low_T15Y13), .B(tie_low_T15Y13), .Y(1025));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10738  (.A(tie_low_T14Y19), .B(tie_low_T14Y19), .Y(1027));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10739  (.A(tie_low_T13Y22), .B(tie_low_T13Y22), .X(1029));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10740  (.A(tie_low_T15Y14), .B(tie_low_T15Y14), .Y(1030));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10741  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(1032));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10742  (.A(tie_low_T13Y22), .B(tie_low_T13Y22), .X(1034));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10743  (.A(tie_low_T15Y14), .B(tie_low_T15Y14), .Y(1035));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10744  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(1037));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10745  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .Y(1038));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10746  (.A(tie_low_T15Y14), .B(tie_low_T15Y14), .Y(1039));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10747  (.A(tie_low_T4Y30), .B(tie_low_T4Y30), .Y(1042));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10748  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .Y(1044));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10749  (.A(1044), .Y(1045));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10750  (.A(tie_low_T7Y31), .B(tie_low_T7Y31), .X(1048));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10751  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1051));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10752  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .X(1053));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10753  (.A(tie_low_T6Y30), .B(tie_low_T6Y30), .Y(1054));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10754  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(1057));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10755  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .X(1059));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10756  (.A(1059), .Y(1060));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10757  (.A(tie_low_T4Y26), .B(tie_low_T4Y26), .X(1063));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10758  (.A(tie_low_T5Y26), .B(tie_low_T5Y26), .Y(1065));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10759  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(1067));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10760  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .X(1068));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10761  (.A(tie_low_T4Y24), .B(tie_low_T4Y24), .Y(1070));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10762  (.A(1070), .Y(1071));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10763  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1074));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10764  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .Y(1075));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10765  (.A(tie_low_T8Y29), .B(tie_low_T8Y29), .X(1077));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10766  (.A(1077), .Y(1078));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10767  (.A(tie_low_T8Y29), .B(tie_low_T8Y29), .Y(1079));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10768  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .X(1080));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10769  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(1081));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10770  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .X(1082));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10771  (.A(tie_low_T8Y29), .B(tie_low_T8Y29), .X(1084));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10772  (.A(tie_low_T6Y31), .B(tie_low_T6Y31), .Y(1086));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10773  (.A(tie_low_T6Y27), .B(tie_low_T6Y27), .X(1089));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10774  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .X(1090));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10775  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1091));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10776  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1092));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10777  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .X(1093));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10778  (.A(tie_low_T6Y26), .B(tie_low_T6Y26), .X(1096));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10779  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .X(1098));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10780  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1099));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10781  (.A(tie_low_T6Y27), .B(tie_low_T6Y27), .Y(1100));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10782  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(1102));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10783  (.A(tie_low_T6Y25), .B(tie_low_T6Y25), .Y(1103));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10784  (.A(tie_low_T4Y28), .B(tie_low_T4Y28), .Y(1104));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10785  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1105));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10786  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .Y(1106));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10787  (.A(1106), .Y(1107));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10788  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .Y(1108));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10789  (.A(tie_low_T6Y27), .B(tie_low_T6Y27), .X(1109));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10790  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .X(1110));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10791  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1111));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10792  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .Y(1112));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10793  (.A(tie_low_T10Y15), .B(tie_low_T10Y15), .Y(1114));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10794  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(1116));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10795  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .X(1117));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10796  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1118));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10797  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(1120));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10798  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(1121));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10799  (.A(1121), .Y(1122));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10800  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1124));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10801  (.A(tie_low_T10Y16), .B(tie_low_T10Y16), .Y(1127));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10802  (.A(1127), .Y(1128));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10803  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1129));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10804  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1131));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10805  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1134));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10806  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(1135));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10807  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(1136));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10808  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1137));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10809  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1138));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10810  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .Y(1139));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10811  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(1140));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10812  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .X(1142));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10813  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(1145));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10814  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1146));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10815  (.A(tie_low_T9Y34), .B(tie_low_T9Y34), .X(1147));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10816  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1148));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10817  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1149));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10818  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1150));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10819  (.A(tie_low_T10Y28), .B(tie_low_T10Y28), .X(1151));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10820  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(1152));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10821  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(1154));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10822  (.A(1154), .Y(1155));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10823  (.A(tie_low_T11Y16), .B(tie_low_T11Y16), .X(1156));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10824  (.A(1156), .Y(1157));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10825  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1158));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10826  (.A(tie_low_T11Y19), .B(tie_low_T11Y19), .X(1159));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10827  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(1162));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10828  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .X(1163));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10829  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .X(1164));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10830  (.A(tie_low_T8Y28), .B(tie_low_T8Y28), .X(1165));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10831  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .X(1166));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10832  (.A(tie_low_T5Y35), .B(tie_low_T5Y35), .X(1167));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10833  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(1168));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10834  (.A(1168), .Y(1169));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10835  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(1170));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10836  (.A(tie_low_T4Y31), .B(tie_low_T4Y31), .X(1171));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10837  (.A(tie_low_T14Y7), .B(tie_low_T14Y7), .Y(1172));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10838  (.A(1172), .Y(1173));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10839  (.A(tie_low_T4Y25), .B(tie_low_T4Y25), .X(1175));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10840  (.A(1175), .Y(1176));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10841  (.A(tie_low_T7Y26), .B(tie_low_T7Y26), .X(1177));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10842  (.A(tie_low_T8Y25), .B(tie_low_T8Y25), .X(1178));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10843  (.A(tie_low_T7Y29), .B(tie_low_T7Y29), .Y(1179));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10844  (.A(tie_low_T8Y23), .B(tie_low_T8Y23), .X(1180));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10845  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1181));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10846  (.A(tie_low_T11Y18), .B(tie_low_T11Y18), .Y(1182));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10847  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .X(1183));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10848  (.A(tie_low_T6Y17), .B(tie_low_T6Y17), .X(1185));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10849  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1186));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10850  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1187));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10851  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(1189));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10852  (.A(1187), .B(1189), .X(1190));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10853  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1191));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10854  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(1192));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10855  (.A(tie_low_T13Y23), .B(tie_low_T13Y23), .X(1194));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10856  (.A(1194), .Y(1195));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10857  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .X(1197));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10858  (.A(640), .B(1197), .X(1198));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10859  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1199));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10860  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1202));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10861  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1203));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10862  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1204));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10863  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(1205));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10864  (.A(629), .B(694), .Y(1206));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10865  (.A(1133), .B(644), .Y(1207));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10866  (.A(1206), .B(1207), .X(1208));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10867  (.A(1205), .B(1208), .X(1209));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10868  (.A(1203), .B(1209), .X(1210));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10869  (.A(1121), .B(1210), .X(1211));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10870  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(1212));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10871  (.A(1212), .Y(1213));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10872  (.A(tie_low_T12Y13), .B(tie_low_T12Y13), .Y(1214));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10873  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1215));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10874  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1217));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10875  (.A(tie_low_T15Y6), .B(tie_low_T15Y6), .Y(1218));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10876  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(1220));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10877  (.A(tie_low_T4Y27), .B(tie_low_T4Y27), .X(1221));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10878  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1222));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10879  (.A(1222), .Y(1223));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10880  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(1224));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10881  (.A(tie_low_T7Y28), .B(tie_low_T7Y28), .X(1225));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10882  (.A(tie_low_T7Y25), .B(tie_low_T7Y25), .X(1226));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10883  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1227));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10884  (.A(tie_low_T19Y33), .B(tie_low_T19Y33), .X(1228));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10885  (.A(1228), .Y(1229));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10886  (.A(tie_low_T17Y2), .B(tie_low_T17Y2), .Y(1231));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10887  (.A(tie_low_T19Y25), .B(tie_low_T19Y25), .X(1233));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10888  (.A(1233), .Y(1234));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10889  (.A(tie_low_T17Y3), .B(tie_low_T17Y3), .Y(1236));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10890  (.A(tie_low_T17Y2), .B(tie_low_T17Y2), .Y(1237));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10891  (.A(tie_low_T18Y13), .B(tie_low_T18Y13), .X(1239));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10892  (.A(tie_low_T16Y10), .B(tie_low_T16Y10), .X(1241));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10893  (.A(tie_low_T19Y25), .B(tie_low_T19Y25), .X(1242));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10894  (.A(tie_low_T14Y14), .B(tie_low_T14Y14), .X(1244));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10895  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(1245));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10896  (.A(tie_low_T16Y7), .B(tie_low_T16Y7), .X(1246));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10897  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .Y(1248));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10898  (.A(tie_low_T17Y1), .B(tie_low_T17Y1), .Y(1250));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10899  (.A(tie_low_T17Y5), .B(tie_low_T17Y5), .Y(1252));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10900  (.A(tie_low_T16Y11), .B(tie_low_T16Y11), .Y(1253));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10901  (.A(tie_low_T17Y9), .B(tie_low_T17Y9), .X(1255));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10902  (.A(tie_low_T16Y15), .B(tie_low_T16Y15), .X(1256));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10903  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .Y(1257));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10904  (.A(tie_low_T16Y20), .B(tie_low_T16Y20), .X(1258));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10905  (.A(tie_low_T15Y28), .B(tie_low_T15Y28), .Y(1260));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10906  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1261));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10907  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(1263));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10908  (.A(1264), .B(1265), .X(1266));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10909  (.A(1266), .Y(1267));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10910  (.A(622), .B(667), .Y(1268));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10911  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1269));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10912  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(1270));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10913  (.A(1266), .B(1270), .X(1271));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10914  (.A(tie_low_T16Y16), .B(tie_low_T16Y16), .Y(1272));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10915  (.A(1272), .Y(1273));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10916  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .Y(1275));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10917  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1277));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10918  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(1278));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10919  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1279));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10920  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1280));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10921  (.A(1280), .Y(1281));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10922  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .Y(1282));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10923  (.A(1271), .B(1282), .X(1283));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10924  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .X(1284));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10925  (.A(1284), .Y(1285));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10926  (.A(tie_low_T12Y13), .B(tie_low_T12Y13), .Y(1286));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10927  (.A(tie_low_T14Y7), .B(tie_low_T14Y7), .X(1287));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10928  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .X(1289));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10929  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1290));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10930  (.A(1290), .Y(1291));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10931  (.A(tie_low_T7Y26), .B(tie_low_T7Y26), .X(1292));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10932  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .X(1293));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10933  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1294));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10934  (.A(tie_low_T6Y16), .B(tie_low_T6Y16), .Y(1296));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10935  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(1297));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10936  (.A(tie_low_T10Y26), .B(tie_low_T10Y26), .X(1298));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10937  (.A(630), .B(1127), .X(1299));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10938  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1300));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10939  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(1301));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10940  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(1303));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10941  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(1304));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10942  (.A(1304), .Y(1305));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10943  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1306));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10944  (.A(1303), .B(1306), .X(1307));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10945  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1308));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10946  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1309));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10947  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(1310));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10948  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(1311));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10949  (.A(1311), .Y(1312));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10950  (.A(tie_low_T11Y15), .B(tie_low_T11Y15), .Y(1313));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10951  (.A(tie_low_T12Y13), .B(tie_low_T12Y13), .X(1314));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10952  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1315));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10953  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1317));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10954  (.A(tie_low_T15Y6), .B(tie_low_T15Y6), .Y(1318));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10955  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(1319));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10956  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1320));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10957  (.A(tie_low_T6Y27), .B(tie_low_T6Y27), .X(1321));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10958  (.A(tie_low_T8Y23), .B(tie_low_T8Y23), .X(1322));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10959  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1323));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10960  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(1324));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10961  (.A(1324), .Y(1325));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10962  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(1326));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10963  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1327));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10964  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1328));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10965  (.A(1130), .B(469), .Y(1329));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10966  (.A(1329), .Y(1330));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10967  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1332));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10968  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1333));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10969  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .X(1334));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10970  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .X(1336));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10971  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(1337));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10972  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(1338));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10973  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1339));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10974  (.A(tie_low_T9Y19), .B(tie_low_T9Y19), .X(1340));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10975  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1341));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10976  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1342));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10977  (.A(1342), .Y(1343));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10978  (.A(tie_low_T12Y13), .B(tie_low_T12Y13), .Y(1344));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10979  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1345));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10980  (.A(tie_low_T14Y7), .B(tie_low_T14Y7), .Y(1347));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10981  (.A(tie_low_T15Y5), .B(tie_low_T15Y5), .Y(1348));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10982  (.A(tie_low_T4Y24), .B(tie_low_T4Y24), .X(1350));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10983  (.A(tie_low_T5Y27), .B(tie_low_T5Y27), .Y(1351));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10984  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .X(1352));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10985  (.A(tie_low_T7Y24), .B(tie_low_T7Y24), .X(1353));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10986  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1354));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10987  (.A(644), .B(1195), .X(1355));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10988  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1356));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10989  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1357));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10990  (.A(1356), .B(1357), .X(1358));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10991  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1360));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10992  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(1361));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10993  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(1362));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10994  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1363));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10995  (.A(1363), .Y(1364));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10996  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(1365));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10997  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .X(1366));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10998  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1367));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$10999  (.A(tie_low_T14Y7), .B(tie_low_T14Y7), .Y(1369));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11000  (.A(tie_low_T15Y5), .B(tie_low_T15Y5), .Y(1370));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11001  (.A(tie_low_T5Y26), .B(tie_low_T5Y26), .Y(1371));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11002  (.A(tie_low_T7Y28), .B(tie_low_T7Y28), .X(1372));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11003  (.A(tie_low_T7Y24), .B(tie_low_T7Y24), .X(1373));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11004  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1374));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11005  (.A(1134), .B(1189), .X(1375));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11006  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1376));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11007  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1377));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11008  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(1378));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11009  (.A(1378), .Y(1379));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11010  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1380));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11011  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(1381));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11012  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(1382));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11013  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(1384));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11014  (.A(tie_low_T15Y5), .B(tie_low_T15Y5), .Y(1385));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11015  (.A(tie_low_T13Y19), .B(tie_low_T13Y19), .X(1388));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11016  (.A(tie_low_T8Y29), .B(tie_low_T8Y29), .X(1390));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11017  (.A(tie_low_T4Y24), .B(tie_low_T4Y24), .X(1391));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11018  (.A(1391), .Y(1392));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11019  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .X(1394));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11020  (.A(tie_low_T6Y27), .B(tie_low_T6Y27), .X(1396));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11021  (.A(tie_low_T7Y29), .B(tie_low_T7Y29), .X(1398));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11022  (.A(tie_low_T8Y28), .B(tie_low_T8Y28), .X(1399));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11023  (.A(tie_low_T7Y29), .B(tie_low_T7Y29), .X(1400));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11024  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .Y(1401));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11025  (.A(tie_low_T8Y29), .B(tie_low_T8Y29), .Y(1402));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11026  (.A(tie_low_T11Y30), .B(tie_low_T11Y30), .X(1403));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11027  (.A(tie_low_T15Y31), .B(tie_low_T15Y31), .X(1405));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11028  (.A(tie_low_T10Y30), .B(tie_low_T10Y30), .X(1407));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11029  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(1408));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11030  (.A(1408), .Y(1409));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11031  (.A(tie_low_T13Y18), .B(tie_low_T13Y18), .X(1411));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11032  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1414));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11033  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1415));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11034  (.A(1415), .Y(1416));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11035  (.A(tie_low_T9Y30), .B(tie_low_T9Y30), .X(1417));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11036  (.A(tie_low_T12Y30), .B(tie_low_T12Y30), .X(1418));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11037  (.A(tie_low_T15Y30), .B(tie_low_T15Y30), .X(1419));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11038  (.A(tie_low_T14Y24), .B(tie_low_T14Y24), .Y(1420));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11039  (.A(1420), .Y(1421));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11040  (.A(tie_low_T15Y30), .B(tie_low_T15Y30), .Y(1423));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11041  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1424));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11042  (.A(tie_low_T5Y36), .B(tie_low_T5Y36), .X(1425));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11043  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1426));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11044  (.A(1426), .Y(1427));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11045  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .Y(1429));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11046  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .X(1430));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11047  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1432));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11048  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(1433));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11049  (.A(1433), .Y(1434));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11050  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .Y(1435));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11051  (.A(tie_low_T5Y33), .B(tie_low_T5Y33), .Y(1437));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11052  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(1439));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11053  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(1440));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11054  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .X(1441));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11055  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .X(1442));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11056  (.A(tie_low_T11Y30), .B(tie_low_T11Y30), .Y(1443));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11057  (.A(1443), .Y(1444));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11058  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(1446));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11059  (.A(1446), .Y(1447));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11060  (.A(tie_low_T7Y29), .B(tie_low_T7Y29), .X(1448));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11061  (.A(tie_low_T13Y19), .B(tie_low_T13Y19), .X(1450));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11062  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .Y(1451));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11063  (.A(1451), .Y(1452));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11064  (.A(tie_low_T13Y18), .B(tie_low_T13Y18), .X(1454));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11065  (.A(tie_low_T4Y31), .B(tie_low_T4Y31), .Y(1457));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11066  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(1458));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11067  (.A(1458), .Y(1459));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11068  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(1461));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11069  (.A(1461), .Y(1462));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11070  (.A(tie_low_T11Y31), .B(tie_low_T11Y31), .Y(1465));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11071  (.A(tie_low_T13Y31), .B(tie_low_T13Y31), .X(1466));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11072  (.A(tie_low_T15Y31), .B(tie_low_T15Y31), .X(1467));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11073  (.A(tie_low_T12Y28), .B(tie_low_T12Y28), .X(1468));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11074  (.A(1468), .Y(1469));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11075  (.A(tie_low_T12Y29), .B(tie_low_T12Y29), .X(1470));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11076  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(1471));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11077  (.A(1471), .Y(1472));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11078  (.A(tie_low_T5Y36), .B(tie_low_T5Y36), .X(1474));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11079  (.A(1474), .Y(1475));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11080  (.A(tie_low_T2Y37), .B(tie_low_T2Y37), .X(1476));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11081  (.A(tie_low_T6Y30), .B(tie_low_T6Y30), .X(1478));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11082  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(1480));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11083  (.A(1480), .Y(1481));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11084  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .Y(1482));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11085  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(1483));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11086  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(1485));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11087  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .X(1486));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11088  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(1487));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11089  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(1489));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11090  (.A(tie_low_T15Y17), .B(tie_low_T15Y17), .Y(1490));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11091  (.A(tie_low_T13Y18), .B(tie_low_T13Y18), .X(1492));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11092  (.A(tie_low_T12Y24), .B(tie_low_T12Y24), .X(1493));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11093  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(1494));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11094  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .Y(1496));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11095  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(1498));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11096  (.A(1498), .Y(1499));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11097  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .X(1500));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11098  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1501));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11099  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(1502));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11100  (.A(1502), .Y(1503));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11101  (.A(tie_low_T13Y18), .B(tie_low_T13Y18), .X(1505));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11102  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1507));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11103  (.A(1507), .Y(1508));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11104  (.A(tie_low_T13Y30), .B(tie_low_T13Y30), .X(1509));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11105  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .X(1510));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11106  (.A(tie_low_T13Y23), .B(tie_low_T13Y23), .Y(1511));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11107  (.A(1511), .Y(1512));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11108  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(1514));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11109  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .X(1515));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11110  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(1516));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11111  (.A(tie_low_T10Y15), .B(tie_low_T10Y15), .X(1518));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11112  (.A(tie_low_T9Y10), .B(tie_low_T9Y10), .X(1519));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11113  (.A(tie_low_T9Y15), .B(tie_low_T9Y15), .X(1520));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11114  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1521));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11115  (.A(1521), .Y(1522));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11116  (.A(tie_low_T16Y11), .B(tie_low_T16Y11), .Y(1524));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11117  (.A(tie_low_T10Y8), .B(tie_low_T10Y8), .X(1526));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11118  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(1527));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11119  (.A(tie_low_T8Y6), .B(tie_low_T8Y6), .X(1528));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11120  (.A(tie_low_T8Y6), .B(tie_low_T8Y6), .Y(1529));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11121  (.A(tie_low_T17Y13), .B(tie_low_T17Y13), .X(1530));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11122  (.A(tie_low_T19Y27), .B(tie_low_T19Y27), .Y(1532));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11123  (.A(tie_low_T17Y18), .B(tie_low_T17Y18), .Y(1533));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11124  (.A(tie_low_T16Y13), .B(tie_low_T16Y13), .X(1534));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11125  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .Y(1535));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11126  (.A(tie_low_T11Y14), .B(tie_low_T11Y14), .Y(1536));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11127  (.A(1536), .Y(1537));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11128  (.A(tie_low_T12Y26), .B(tie_low_T12Y26), .Y(1538));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11129  (.A(1538), .Y(1539));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11130  (.A(607), .B(667), .Y(1540));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11131  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1541));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11132  (.A(1139), .B(1541), .X(1542));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11133  (.A(tie_low_T15Y13), .B(tie_low_T15Y13), .X(1544));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11134  (.A(tie_low_T12Y10), .B(tie_low_T12Y10), .Y(1545));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11135  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(1546));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11136  (.A(tie_low_T16Y13), .B(tie_low_T16Y13), .X(1547));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11137  (.A(tie_low_T15Y15), .B(tie_low_T15Y15), .Y(1548));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11138  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(1549));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11139  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(1550));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11140  (.A(1542), .B(1550), .X(1551));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11141  (.A(1539), .B(1551), .X(1552));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11142  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(1553));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11143  (.A(tie_low_T8Y16), .B(tie_low_T8Y16), .X(1554));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11144  (.A(tie_low_T12Y13), .B(tie_low_T12Y13), .Y(1556));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11145  (.A(tie_low_T10Y11), .B(tie_low_T10Y11), .Y(1557));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11146  (.A(1557), .Y(1558));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11147  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .X(1559));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11148  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(1560));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11149  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .X(1561));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11150  (.A(tie_low_T8Y36), .B(tie_low_T8Y36), .X(1562));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11151  (.A(1563), .B(1303), .X(1564));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11152  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(1566));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11153  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .X(1567));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11154  (.A(tie_low_T10Y10), .B(tie_low_T10Y10), .X(1568));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11155  (.A(1568), .Y(1569));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11156  (.A(tie_low_T10Y26), .B(tie_low_T10Y26), .X(1570));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11157  (.A(1570), .Y(1571));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11158  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .X(1572));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11159  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1573));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11160  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .X(1574));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11161  (.A(626), .B(1574), .X(1575));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11162  (.A(tie_low_T11Y16), .B(tie_low_T11Y16), .X(1576));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11163  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(1577));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11164  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .X(1579));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11165  (.A(1576), .B(1579), .X(1580));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11166  (.A(1575), .B(1580), .X(1581));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11167  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .X(1582));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11168  (.A(1582), .Y(1583));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11169  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(1584));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11170  (.A(tie_low_T7Y11), .B(tie_low_T7Y11), .X(1585));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11171  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .Y(1586));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11172  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .Y(1587));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11173  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .Y(1588));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11174  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(1589));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11175  (.A(1589), .Y(1590));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11176  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(1591));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11177  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1592));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11178  (.A(1592), .Y(1593));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11179  (.A(tie_low_T3Y37), .B(tie_low_T3Y37), .Y(1594));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11180  (.A(tie_low_T12Y11), .B(tie_low_T12Y11), .Y(1595));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11181  (.A(1595), .Y(1596));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11182  (.A(tie_low_T12Y11), .B(tie_low_T12Y11), .Y(1597));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11183  (.A(1597), .Y(1598));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11184  (.A(1599), .B(1187), .X(1600));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11185  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .X(1601));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11186  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .X(1602));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11187  (.A(tie_low_T17Y28), .B(tie_low_T17Y28), .X(1603));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11188  (.A(tie_low_T13Y21), .B(tie_low_T13Y21), .X(1604));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11189  (.A(1604), .Y(1605));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11190  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1606));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11191  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1607));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11192  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1608));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11193  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1609));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11194  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .Y(1610));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11195  (.A(620), .B(1610), .X(1611));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11196  (.A(tie_low_T10Y18), .B(tie_low_T10Y18), .X(1612));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11197  (.A(1611), .B(1612), .X(1613));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11198  (.A(1297), .B(1564), .X(1614));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11199  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .X(1615));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11200  (.A(tie_low_T13Y24), .B(tie_low_T13Y24), .X(1616));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11201  (.A(1616), .Y(1617));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11202  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .Y(1618));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11203  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(1619));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11204  (.A(tie_low_T12Y22), .B(tie_low_T12Y22), .Y(1620));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11205  (.A(1620), .Y(1621));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11206  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(1622));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11207  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1623));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11208  (.A(tie_low_T8Y26), .B(tie_low_T8Y26), .Y(1624));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11209  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(1625));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11210  (.A(tie_low_T3Y37), .B(tie_low_T3Y37), .X(1626));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11211  (.A(1626), .Y(1627));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11212  (.A(tie_low_T4Y32), .B(tie_low_T4Y32), .Y(1628));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11213  (.A(tie_low_T7Y18), .B(tie_low_T7Y18), .Y(1629));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11214  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(1630));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11215  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1631));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11216  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1632));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11217  (.A(tie_low_T12Y10), .B(tie_low_T12Y10), .Y(1633));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11218  (.A(tie_low_T11Y15), .B(tie_low_T11Y15), .Y(1634));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11219  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(1635));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11220  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .Y(1636));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11221  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(1637));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11222  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1638));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11223  (.A(1638), .Y(1639));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11224  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1640));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11225  (.A(1634), .B(1638), .X(1641));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11226  (.A(1620), .B(1641), .Y(1642));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11227  (.A(tie_low_T10Y16), .B(tie_low_T10Y16), .X(1643));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11228  (.A(1621), .B(1643), .Y(1644));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11229  (.A(1642), .B(1644), .Y(1645));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11230  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1646));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11231  (.A(tie_low_T11Y15), .B(tie_low_T11Y15), .X(1647));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11232  (.A(1647), .Y(1648));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11233  (.A(tie_low_T11Y16), .B(tie_low_T11Y16), .Y(1649));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11234  (.A(1649), .Y(1650));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11235  (.A(tie_low_T14Y34), .B(tie_low_T14Y34), .Y(1651));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11236  (.A(tie_low_T21Y70), .B(tie_low_T21Y70), .X(1652));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11237  (.A(tie_low_T20Y45), .B(tie_low_T20Y45), .Y(1653));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11238  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(1654));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11239  (.A(tie_low_T13Y22), .B(tie_low_T13Y22), .X(1655));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11240  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(1656));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11241  (.A(tie_low_T12Y22), .B(tie_low_T12Y22), .Y(1657));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11242  (.A(1657), .Y(1658));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11243  (.A(1643), .B(1657), .X(1659));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11244  (.A(1641), .B(1658), .X(1660));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11245  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1661));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11246  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1662));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11247  (.A(tie_low_T10Y26), .B(tie_low_T10Y26), .X(1663));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11248  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(1664));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11249  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(1665));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11250  (.A(401), .B(1665), .Y(1666));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11251  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .Y(1667));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11252  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1668));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11253  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1669));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11254  (.A(1669), .Y(1670));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11255  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .Y(1671));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11256  (.A(1671), .Y(1672));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11257  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1673));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11258  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(1674));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11259  (.A(1674), .Y(1675));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11260  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1676));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11261  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(1677));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11262  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1678));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11263  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1679));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11264  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(1680));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11265  (.A(tie_low_T7Y18), .B(tie_low_T7Y18), .Y(1681));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11266  (.A(tie_low_T7Y23), .B(tie_low_T7Y23), .X(1682));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11267  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1683));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11268  (.A(tie_low_T5Y33), .B(tie_low_T5Y33), .Y(1684));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11269  (.A(tie_low_T13Y22), .B(tie_low_T13Y22), .X(1685));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11270  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(1686));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11271  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(1687));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11272  (.A(1687), .Y(1688));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11273  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(1689));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11274  (.A(1643), .B(1688), .Y(1690));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11275  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(1691));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11276  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1692));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11277  (.A(1692), .Y(1693));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11278  (.A(tie_low_T11Y29), .B(tie_low_T11Y29), .X(1694));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11279  (.A(191), .B(1575), .Y(1695));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11280  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(1696));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11281  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(1697));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11282  (.A(1697), .Y(1698));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11283  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(1699));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11284  (.A(1586), .B(1699), .X(1700));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11285  (.A(1700), .Y(1701));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11286  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(1702));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11287  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1703));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11288  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1704));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11289  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1705));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11290  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1706));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11291  (.A(tie_low_T8Y23), .B(tie_low_T8Y23), .X(1707));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11292  (.A(tie_low_T8Y23), .B(tie_low_T8Y23), .Y(1708));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11293  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(1709));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11294  (.A(tie_low_T7Y21), .B(tie_low_T7Y21), .X(1710));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11295  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .X(1711));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11296  (.A(tie_low_T9Y19), .B(tie_low_T9Y19), .Y(1712));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11297  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1713));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11298  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .Y(1714));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11299  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(1715));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11300  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(1716));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11301  (.A(1716), .Y(1717));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11302  (.A(1643), .B(1716), .X(1718));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11303  (.A(1641), .B(1717), .X(1719));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11304  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1720));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11305  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1721));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11306  (.A(tie_low_T11Y30), .B(tie_low_T11Y30), .X(1722));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11307  (.A(169), .B(1575), .Y(1723));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11308  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .Y(1724));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11309  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(1725));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11310  (.A(1725), .Y(1726));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11311  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(1727));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11312  (.A(1586), .B(1727), .X(1728));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11313  (.A(1728), .Y(1729));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11314  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(1730));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11315  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1731));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11316  (.A(1731), .Y(1732));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11317  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(1733));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11318  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1734));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11319  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1735));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11320  (.A(1735), .Y(1736));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11321  (.A(tie_low_T8Y20), .B(tie_low_T8Y20), .Y(1737));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11322  (.A(tie_low_T8Y20), .B(tie_low_T8Y20), .X(1738));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11323  (.A(1738), .Y(1739));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11324  (.A(tie_low_T7Y20), .B(tie_low_T7Y20), .Y(1740));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11325  (.A(tie_low_T7Y18), .B(tie_low_T7Y18), .Y(1741));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11326  (.A(tie_low_T8Y19), .B(tie_low_T8Y19), .X(1742));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11327  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1743));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11328  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1744));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11329  (.A(tie_low_T13Y24), .B(tie_low_T13Y24), .X(1745));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11330  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(1746));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11331  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(1747));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11332  (.A(1747), .Y(1748));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11333  (.A(1641), .B(1747), .Y(1749));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11334  (.A(1643), .B(1748), .Y(1750));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11335  (.A(1749), .B(1750), .Y(1751));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11336  (.A(tie_low_T11Y16), .B(tie_low_T11Y16), .Y(1752));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11337  (.A(1752), .Y(1753));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11338  (.A(tie_low_T10Y28), .B(tie_low_T10Y28), .X(1754));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11339  (.A(145), .B(1575), .Y(1755));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11340  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(1756));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11341  (.A(334), .B(1756), .Y(1757));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11342  (.A(1757), .Y(1758));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11343  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(1759));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11344  (.A(1586), .B(1759), .X(1760));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11345  (.A(1760), .Y(1761));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11346  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .Y(1762));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11347  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1763));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11348  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1764));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11349  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(1765));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11350  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1766));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11351  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1767));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11352  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1768));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11353  (.A(tie_low_T8Y20), .B(tie_low_T8Y20), .Y(1769));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11354  (.A(tie_low_T7Y20), .B(tie_low_T7Y20), .X(1770));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11355  (.A(tie_low_T7Y18), .B(tie_low_T7Y18), .X(1771));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11356  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .Y(1772));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11357  (.A(1753), .B(1772), .X(1773));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11358  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1774));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11359  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1775));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11360  (.A(1775), .Y(1776));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11361  (.A(tie_low_T13Y24), .B(tie_low_T13Y24), .X(1777));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11362  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(1778));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11363  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .Y(1779));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11364  (.A(1779), .Y(1780));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11365  (.A(1641), .B(1779), .Y(1781));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11366  (.A(1643), .B(1780), .Y(1782));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11367  (.A(1781), .B(1782), .Y(1783));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11368  (.A(tie_low_T11Y16), .B(tie_low_T11Y16), .Y(1784));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11369  (.A(1784), .Y(1785));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11370  (.A(tie_low_T10Y29), .B(tie_low_T10Y29), .X(1786));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11371  (.A(518), .B(1575), .Y(1787));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11372  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(1788));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11373  (.A(tie_low_T10Y16), .B(tie_low_T10Y16), .Y(1789));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11374  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(1790));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11375  (.A(1790), .Y(1791));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11376  (.A(tie_low_T9Y23), .B(tie_low_T9Y23), .Y(1792));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11377  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1793));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11378  (.A(1793), .Y(1794));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11379  (.A(tie_low_T9Y23), .B(tie_low_T9Y23), .Y(1795));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11380  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1796));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11381  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1797));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11382  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(1798));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11383  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1799));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11384  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .X(1800));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11385  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .Y(1801));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11386  (.A(tie_low_T8Y21), .B(tie_low_T8Y21), .Y(1802));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11387  (.A(tie_low_T7Y21), .B(tie_low_T7Y21), .X(1803));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11388  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .X(1804));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11389  (.A(tie_low_T9Y19), .B(tie_low_T9Y19), .Y(1805));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11390  (.A(1785), .B(1805), .X(1806));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11391  (.A(tie_low_T13Y23), .B(tie_low_T13Y23), .X(1807));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11392  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(1808));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11393  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(1809));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11394  (.A(1809), .Y(1810));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11395  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(1811));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11396  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .X(1812));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11397  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(1813));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11398  (.A(tie_low_T7Y24), .B(tie_low_T7Y24), .X(1814));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11399  (.A(tie_low_T10Y29), .B(tie_low_T10Y29), .X(1815));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11400  (.A(286), .B(1575), .Y(1816));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11401  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(1817));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11402  (.A(tie_low_T11Y20), .B(tie_low_T11Y20), .Y(1818));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11403  (.A(tie_low_T10Y16), .B(tie_low_T10Y16), .Y(1819));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11404  (.A(1819), .Y(1820));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11405  (.A(tie_low_T9Y27), .B(tie_low_T9Y27), .Y(1821));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11406  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .X(1822));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11407  (.A(1822), .Y(1823));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11408  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(1824));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11409  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .X(1825));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11410  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1826));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11411  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1827));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11412  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1828));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11413  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(1829));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11414  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .X(1830));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11415  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1831));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11416  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .Y(1832));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11417  (.A(tie_low_T7Y21), .B(tie_low_T7Y21), .Y(1833));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11418  (.A(tie_low_T7Y19), .B(tie_low_T7Y19), .Y(1834));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11419  (.A(tie_low_T4Y32), .B(tie_low_T4Y32), .Y(1835));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11420  (.A(tie_low_T13Y23), .B(tie_low_T13Y23), .X(1836));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11421  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(1837));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11422  (.A(tie_low_T12Y22), .B(tie_low_T12Y22), .Y(1838));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11423  (.A(1838), .Y(1839));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11424  (.A(1643), .B(1838), .X(1840));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11425  (.A(1641), .B(1839), .X(1841));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11426  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .Y(1842));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11427  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1843));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11428  (.A(tie_low_T7Y21), .B(tie_low_T7Y21), .Y(1844));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11429  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(1845));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11430  (.A(516), .B(1575), .Y(1846));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11431  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .Y(1847));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11432  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(1848));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11433  (.A(1848), .Y(1849));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11434  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(1850));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11435  (.A(1586), .B(1850), .X(1851));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11436  (.A(1851), .Y(1852));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11437  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1853));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11438  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1854));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11439  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(1855));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11440  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1856));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11441  (.A(tie_low_T10Y21), .B(tie_low_T10Y21), .Y(1857));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11442  (.A(tie_low_T8Y19), .B(tie_low_T8Y19), .X(1858));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11443  (.A(tie_low_T8Y19), .B(tie_low_T8Y19), .Y(1859));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11444  (.A(tie_low_T8Y19), .B(tie_low_T8Y19), .Y(1860));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11445  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .Y(1861));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11446  (.A(tie_low_T7Y19), .B(tie_low_T7Y19), .Y(1862));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11447  (.A(tie_low_T8Y20), .B(tie_low_T8Y20), .Y(1863));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11448  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(1864));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11449  (.A(tie_low_T7Y24), .B(tie_low_T7Y24), .Y(1865));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11450  (.A(tie_low_T10Y16), .B(tie_low_T10Y16), .Y(1866));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11451  (.A(tie_low_T8Y15), .B(tie_low_T8Y15), .Y(1867));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11452  (.A(tie_low_T8Y15), .B(tie_low_T8Y15), .X(1868));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11453  (.A(tie_low_T9Y10), .B(tie_low_T9Y10), .Y(1869));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11454  (.A(tie_low_T8Y12), .B(tie_low_T8Y12), .Y(1870));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11455  (.A(tie_low_T7Y23), .B(tie_low_T7Y23), .X(1871));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11456  (.A(tie_low_T4Y33), .B(tie_low_T4Y33), .Y(1872));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11457  (.A(tie_low_T6Y25), .B(tie_low_T6Y25), .X(1873));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11458  (.A(tie_low_T4Y34), .B(tie_low_T4Y34), .Y(1874));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11459  (.A(1874), .Y(1875));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11460  (.A(tie_low_T0Y46), .B(tie_low_T0Y46), .Y(1876));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11461  (.A(tie_low_T1Y45), .B(tie_low_T1Y45), .Y(1877));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11462  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1878));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11463  (.A(tie_low_T8Y23), .B(tie_low_T8Y23), .Y(1879));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11464  (.A(1879), .Y(1880));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11465  (.A(tie_low_T2Y41), .B(tie_low_T2Y41), .Y(1881));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11466  (.A(tie_low_T5Y33), .B(tie_low_T5Y33), .Y(1882));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11467  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .Y(1883));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11468  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1884));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11469  (.A(tie_low_T5Y33), .B(tie_low_T5Y33), .Y(1885));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11470  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(1887));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11471  (.A(1887), .Y(1888));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11472  (.A(tie_low_T1Y45), .B(tie_low_T1Y45), .X(1889));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11473  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(1890));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11474  (.A(tie_low_T1Y43), .B(tie_low_T1Y43), .X(1891));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11475  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(1892));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11476  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(1893));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11477  (.A(tie_low_T0Y47), .B(tie_low_T0Y47), .Y(1894));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11478  (.A(tie_low_T2Y42), .B(tie_low_T2Y42), .X(1895));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11479  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(1896));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11480  (.A(1896), .Y(1897));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11481  (.A(tie_low_T1Y44), .B(tie_low_T1Y44), .Y(1898));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11482  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1899));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11483  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .Y(1900));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11484  (.A(1900), .Y(1901));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11485  (.A(tie_low_T3Y40), .B(tie_low_T3Y40), .Y(1902));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11486  (.A(tie_low_T6Y31), .B(tie_low_T6Y31), .Y(1903));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11487  (.A(1691), .B(1712), .Y(1904));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11488  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .Y(1905));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11489  (.A(1905), .Y(1906));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11490  (.A(tie_low_T2Y42), .B(tie_low_T2Y42), .Y(1907));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11491  (.A(tie_low_T5Y35), .B(tie_low_T5Y35), .Y(1908));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11492  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .X(1909));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11493  (.A(tie_low_T5Y35), .B(tie_low_T5Y35), .Y(1910));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11494  (.A(1910), .Y(1911));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11495  (.A(tie_low_T2Y42), .B(tie_low_T2Y42), .Y(1912));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11496  (.A(tie_low_T1Y46), .B(tie_low_T1Y46), .Y(1913));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11497  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .X(1914));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11498  (.A(1914), .Y(1915));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11499  (.A(tie_low_T13Y26), .B(tie_low_T13Y26), .Y(1916));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11500  (.A(tie_low_T7Y36), .B(tie_low_T7Y36), .Y(1917));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11501  (.A(tie_low_T7Y36), .B(tie_low_T7Y36), .X(1918));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11502  (.A(tie_low_T11Y47), .B(tie_low_T11Y47), .Y(1919));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11503  (.A(tie_low_T21Y70), .B(tie_low_T21Y70), .X(1920));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11504  (.A(tie_low_T10Y60), .B(tie_low_T10Y60), .Y(1921));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11505  (.A(1921), .Y(1922));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11506  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(1924));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11507  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(1925));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11508  (.A(tie_low_T13Y39), .B(tie_low_T13Y39), .Y(1926));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11509  (.A(tie_low_T7Y20), .B(tie_low_T7Y20), .Y(1927));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11510  (.A(tie_low_T4Y32), .B(tie_low_T4Y32), .Y(1928));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11511  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(1929));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11512  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .X(1930));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11513  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(1931));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11514  (.A(1931), .Y(1932));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11515  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(1933));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11516  (.A(tie_low_T0Y49), .B(tie_low_T0Y49), .Y(1934));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11517  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(1935));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11518  (.A(1935), .Y(1936));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11519  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(1937));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11520  (.A(39), .B(1890), .Y(1938));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11521  (.A(1937), .B(1938), .Y(1939));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11522  (.A(1939), .Y(1940));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11523  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(1941));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11524  (.A(39), .B(1885), .Y(1942));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11525  (.A(1941), .B(1942), .Y(1943));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11526  (.A(1943), .Y(1944));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11527  (.A(tie_low_T1Y43), .B(tie_low_T1Y43), .X(1945));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11528  (.A(tie_low_T3Y41), .B(tie_low_T3Y41), .Y(1946));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11529  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .Y(1947));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11530  (.A(39), .B(169), .X(1948));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11531  (.A(1947), .B(1948), .Y(1949));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11532  (.A(1949), .Y(1950));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11533  (.A(tie_low_T2Y41), .B(tie_low_T2Y41), .X(1951));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11534  (.A(1907), .B(1951), .Y(1952));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11535  (.A(39), .B(191), .X(1953));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11536  (.A(39), .B(1952), .Y(1954));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11537  (.A(1953), .B(1954), .Y(1955));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11538  (.A(1955), .Y(1956));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11539  (.A(tie_low_T2Y42), .B(tie_low_T2Y42), .X(1957));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11540  (.A(1912), .B(1957), .Y(1958));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11541  (.A(39), .B(213), .X(1959));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11542  (.A(39), .B(1958), .Y(1960));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11543  (.A(1959), .B(1960), .Y(1961));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11544  (.A(1961), .Y(1962));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11545  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(1964));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11546  (.A(39), .B(1594), .Y(1965));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11547  (.A(tie_low_T13Y39), .B(tie_low_T13Y39), .Y(1966));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11548  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(1967));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11549  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .X(1968));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11550  (.A(tie_low_T9Y10), .B(tie_low_T9Y10), .Y(1969));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11551  (.A(tie_low_T8Y14), .B(tie_low_T8Y14), .Y(1970));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11552  (.A(tie_low_T7Y36), .B(tie_low_T7Y36), .X(1971));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11553  (.A(tie_low_T13Y26), .B(tie_low_T13Y26), .Y(1972));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11554  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .X(1973));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11555  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1974));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11556  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1975));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11557  (.A(1952), .B(1958), .Y(1976));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11558  (.A(1888), .B(1976), .Y(1977));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11559  (.A(39), .B(1977), .Y(1978));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11560  (.A(tie_low_T10Y59), .B(tie_low_T10Y59), .Y(1979));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11561  (.A(tie_low_T10Y40), .B(tie_low_T10Y40), .Y(1980));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11562  (.A(tie_low_T5Y45), .B(tie_low_T5Y45), .Y(1981));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11563  (.A(1981), .Y(1982));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11564  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(1984));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11565  (.A(tie_low_T0Y40), .B(tie_low_T0Y40), .Y(1986));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11566  (.A(tie_low_T17Y36), .B(tie_low_T17Y36), .X(1987));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11567  (.A(tie_low_T8Y24), .B(tie_low_T8Y24), .Y(1989));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11568  (.A(tie_low_T13Y30), .B(tie_low_T13Y30), .Y(1990));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11569  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(1991));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11570  (.A(1991), .Y(1992));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11571  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .X(1993));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11572  (.A(1993), .Y(1994));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11573  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(1996));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11574  (.A(tie_low_T18Y0), .B(tie_low_T18Y0), .Y(1997));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11575  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .X(1998));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11576  (.A(tie_low_T14Y32), .B(tie_low_T14Y32), .Y(1999));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11577  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .X(2001));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11578  (.A(tie_low_T8Y27), .B(tie_low_T8Y27), .Y(2002));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11579  (.A(tie_low_T15Y38), .B(tie_low_T15Y38), .Y(2003));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11580  (.A(tie_low_T13Y29), .B(tie_low_T13Y29), .Y(2004));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11581  (.A(tie_low_T15Y22), .B(tie_low_T15Y22), .Y(2005));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11582  (.A(tie_low_T15Y16), .B(tie_low_T15Y16), .Y(2006));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11583  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .X(2007));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11584  (.A(2007), .Y(2008));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11585  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .Y(2010));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11586  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .X(2011));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11587  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(2012));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11588  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .Y(2013));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11589  (.A(tie_low_T35Y60), .B(tie_low_T35Y60), .Y(2015));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11590  (.A(tie_low_T14Y8), .B(tie_low_T14Y8), .Y(2017));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11591  (.A(tie_low_T19Y26), .B(tie_low_T19Y26), .Y(2018));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11592  (.A(tie_low_T8Y9), .B(tie_low_T8Y9), .Y(2020));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11593  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(2022));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11594  (.A(tie_low_T5Y10), .B(tie_low_T5Y10), .Y(2023));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11595  (.A(661), .B(2023), .Y(2024));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11596  (.A(2013), .B(2024), .Y(2025));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11597  (.A(469), .B(2025), .Y(2026));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11598  (.A(1015), .B(469), .X(2027));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11599  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(2028));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11600  (.A(2028), .Y(2029));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11601  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2030));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11602  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(2031));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11603  (.A(tie_low_T14Y16), .B(tie_low_T14Y16), .Y(2032));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11604  (.A(tie_low_T9Y19), .B(tie_low_T9Y19), .X(2033));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11605  (.A(2033), .Y(2034));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11606  (.A(tie_low_T9Y10), .B(tie_low_T9Y10), .X(2035));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11607  (.A(tie_low_T7Y15), .B(tie_low_T7Y15), .Y(2036));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11608  (.A(tie_low_T0Y20), .B(tie_low_T0Y20), .X(116));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11609  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .Y(2037));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11610  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .X(2040));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11611  (.A(150), .B(2040), .Y(2041));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11612  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(2042));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11613  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .X(2044));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11614  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(2045));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11615  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(2046));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11616  (.A(tie_low_T13Y18), .B(tie_low_T13Y18), .Y(2047));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11617  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(2048));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11618  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2049));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11619  (.A(tie_low_T13Y41), .B(tie_low_T13Y41), .Y(2050));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11620  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .Y(2051));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11621  (.A(2051), .Y(2052));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11622  (.A(tie_low_T12Y56), .B(tie_low_T12Y56), .Y(2053));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11623  (.A(tie_low_T15Y89), .B(tie_low_T15Y89), .X(108));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11624  (.A(tie_low_T11Y43), .B(tie_low_T11Y43), .X(2054));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11625  (.A(286), .B(2045), .Y(2055));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11626  (.A(2055), .Y(2056));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11627  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2057));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11628  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(2058));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11629  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2059));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11630  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2060));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11631  (.A(2060), .Y(2061));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11632  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2062));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11633  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2063));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11634  (.A(2063), .Y(2064));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11635  (.A(tie_low_T19Y89), .B(tie_low_T19Y89), .Y(109));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11636  (.A(tie_low_T12Y43), .B(tie_low_T12Y43), .X(2065));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11637  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2066));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11638  (.A(2066), .Y(2067));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11639  (.A(518), .B(2045), .Y(2068));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11640  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2069));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11641  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(2070));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11642  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2071));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11643  (.A(2071), .Y(2072));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11644  (.A(2068), .B(2072), .Y(2073));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11645  (.A(2067), .B(2073), .X(2074));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11646  (.A(2074), .Y(2075));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11647  (.A(tie_low_T23Y89), .B(tie_low_T23Y89), .Y(110));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11648  (.A(tie_low_T9Y34), .B(tie_low_T9Y34), .X(2076));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11649  (.A(145), .B(2045), .Y(2077));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11650  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2078));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11651  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(2079));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11652  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2080));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11653  (.A(tie_low_T17Y41), .B(tie_low_T17Y41), .Y(2081));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11654  (.A(tie_low_T10Y24), .B(tie_low_T10Y24), .Y(2082));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11655  (.A(2082), .Y(2083));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11656  (.A(tie_low_T18Y61), .B(tie_low_T18Y61), .Y(2084));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11657  (.A(tie_low_T27Y89), .B(tie_low_T27Y89), .X(111));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11658  (.A(tie_low_T13Y43), .B(tie_low_T13Y43), .X(2085));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11659  (.A(169), .B(2045), .Y(2086));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11660  (.A(2086), .Y(2087));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11661  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(2088));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11662  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2089));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11663  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2090));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11664  (.A(tie_low_T17Y29), .B(tie_low_T17Y29), .X(2091));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11665  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(2093));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11666  (.A(tie_low_T12Y22), .B(tie_low_T12Y22), .Y(2094));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11667  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .X(2095));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11668  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .X(2096));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11669  (.A(2096), .Y(2097));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11670  (.A(tie_low_T31Y89), .B(tie_low_T31Y89), .Y(112));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11671  (.A(tie_low_T14Y43), .B(tie_low_T14Y43), .X(2098));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11672  (.A(191), .B(2045), .Y(2099));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11673  (.A(2099), .Y(2100));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11674  (.A(150), .B(2091), .Y(2101));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11675  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2102));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11676  (.A(tie_low_T12Y23), .B(tie_low_T12Y23), .Y(2103));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11677  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2104));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11678  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(2105));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11679  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(2106));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11680  (.A(2106), .Y(2107));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11681  (.A(tie_low_T35Y89), .B(tie_low_T35Y89), .Y(113));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11682  (.A(tie_low_T8Y30), .B(tie_low_T8Y30), .X(2108));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11683  (.A(213), .B(2045), .Y(2109));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11684  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2111));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11685  (.A(2111), .Y(2112));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11686  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2113));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11687  (.A(2113), .Y(2114));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11688  (.A(tie_low_T12Y24), .B(tie_low_T12Y24), .Y(2115));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11689  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .Y(2116));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11690  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .X(2117));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11691  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .X(2118));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11692  (.A(2118), .Y(2119));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11693  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(114));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11694  (.A(tie_low_T8Y31), .B(tie_low_T8Y31), .X(2120));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11695  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2122));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11696  (.A(2122), .Y(2123));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11697  (.A(tie_low_T9Y23), .B(tie_low_T9Y23), .X(2124));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11698  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(2125));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11699  (.A(tie_low_T14Y25), .B(tie_low_T14Y25), .Y(2126));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11700  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .Y(2127));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11701  (.A(tie_low_T12Y24), .B(tie_low_T12Y24), .Y(2128));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11702  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .X(2129));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11703  (.A(tie_low_T11Y23), .B(tie_low_T11Y23), .X(2130));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11704  (.A(2130), .Y(2131));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11705  (.A(tie_low_T0Y10), .B(tie_low_T0Y10), .Y(115));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11706  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .Y(2132));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$11707  (.A(2132), .Y(2133));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9277  (.A(2134), .Y(705));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9278  (.A(2135), .Y(595));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9279  (.A(2136), .Y(587));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9280  (.A(2110), .Y(1254));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9281  (.A(1988), .Y(1983));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9282  (.A(60), .Y(1531));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9283  (.A(462), .Y(2137));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9284  (.A(2043), .Y(2038));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9285  (.A(453), .Y(459));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9286  (.A(2021), .Y(2019));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9287  (.A(2014), .Y(2016));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9288  (.A(2138), .Y(2139));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9289  (.A(544), .Y(484));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9290  (.A(39), .Y(433));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9291  (.A(448), .Y(1259));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9292  (.A(2121), .Y(496));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9293  (.A(531), .Y(1240));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9294  (.A(577), .Y(1243));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9295  (.A(1006), .Y(2140));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9296  (.A(1010), .Y(2141));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9297  (.A(1013), .Y(2142));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9298  (.A(1019), .Y(2143));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9299  (.A(1023), .Y(2144));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9300  (.A(1031), .Y(2145));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9301  (.A(1036), .Y(2146));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9302  (.A(2147), .Y(1422));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9303  (.A(234), .Y(236));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9304  (.A(516), .Y(263));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9305  (.A(518), .Y(309));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9306  (.A(169), .Y(171));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9307  (.A(213), .Y(215));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9308  (.A(44), .Y(456));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9309  (.A(3), .Y(1002));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9310  (.A(2148), .Y(1247));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9311  (.A(tie_low_T13Y11), .B(tie_low_T13Y11), .X(488));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9312  (.A(488), .Y(690));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9313  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(2151));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9314  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(608));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9315  (.A(2151), .B(608), .X(666));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9316  (.A(488), .B(666), .X(2039));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9317  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(2153));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9318  (.A(2151), .B(2153), .X(2154));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9319  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .X(614));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9320  (.A(614), .Y(1123));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9321  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .X(1274));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9322  (.A(1274), .Y(2156));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9323  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(1599));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9324  (.A(tie_low_T12Y10), .B(tie_low_T12Y10), .X(605));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9325  (.A(605), .Y(2157));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9326  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(641));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9327  (.A(2153), .B(641), .X(1153));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9328  (.A(tie_low_T9Y19), .B(tie_low_T9Y19), .X(1160));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9329  (.A(488), .B(2154), .X(1161));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9330  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(609));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9331  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(642));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9332  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(654));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9333  (.A(488), .B(654), .X(1132));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9334  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(1264));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9335  (.A(2039), .B(1160), .Y(1563));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9336  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(2160));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9337  (.A(1563), .B(2160), .X(603));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9338  (.A(603), .Y(719));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9339  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(2161));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9340  (.A(tie_low_T11Y17), .B(tie_low_T11Y17), .X(623));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9341  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(1125));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9342  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .X(2162));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9343  (.A(641), .B(2162), .X(2163));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9344  (.A(488), .B(2163), .X(629));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9345  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .Y(2164));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9346  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(606));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9347  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2165));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9348  (.A(2165), .Y(697));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9349  (.A(488), .B(1153), .X(1188));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9350  (.A(2165), .B(1188), .Y(634));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9351  (.A(2151), .B(2162), .X(489));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9352  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(694));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9353  (.A(694), .Y(1265));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9354  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .X(1302));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9355  (.A(694), .B(1302), .Y(2166));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9356  (.A(2164), .B(2166), .X(2167));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9357  (.A(634), .B(2167), .X(2168));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9358  (.A(603), .B(2168), .X(2169));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9359  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(1066));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9360  (.A(1066), .Y(472));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9361  (.A(2169), .B(472), .X(2170));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9362  (.A(608), .B(641), .X(615));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9363  (.A(tie_low_T15Y8), .B(tie_low_T15Y8), .X(611));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9364  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .X(1133));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9365  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(639));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9366  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(617));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9367  (.A(1133), .B(617), .Y(1359));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9368  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(1130));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9369  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(2171));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9370  (.A(1130), .B(2171), .Y(1276));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9371  (.A(1359), .B(1276), .X(1565));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9372  (.A(1565), .Y(2172));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9373  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(2173));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9374  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .X(2174));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9375  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .Y(2176));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9376  (.A(tie_low_T11Y15), .B(tie_low_T11Y15), .Y(2177));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9377  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2178));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9378  (.A(2169), .B(2178), .X(2179));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9379  (.A(2179), .Y(2180));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9380  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(588));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9381  (.A(588), .Y(737));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9382  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(1335));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9383  (.A(1335), .Y(1200));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9384  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(1143));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9385  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2182));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9386  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(2183));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9387  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(2184));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9388  (.A(tie_low_T6Y15), .B(tie_low_T6Y15), .Y(2185));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9389  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .X(2186));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9390  (.A(tie_low_T7Y28), .B(tie_low_T7Y28), .X(2187));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9391  (.A(39), .B(2187), .Y(2188));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9392  (.A(2188), .Y(2189));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9393  (.A(tie_low_T13Y20), .B(tie_low_T13Y20), .X(2190));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9394  (.A(tie_low_T11Y15), .B(tie_low_T11Y15), .Y(2191));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9395  (.A(tie_low_T12Y14), .B(tie_low_T12Y14), .Y(2192));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9396  (.A(2192), .Y(2193));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9397  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(600));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9398  (.A(600), .Y(593));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9399  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2194));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9400  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .X(2195));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9401  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .X(2198));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9402  (.A(tie_low_T12Y17), .B(tie_low_T12Y17), .X(2200));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9403  (.A(tie_low_T15Y14), .B(tie_low_T15Y14), .X(2201));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9404  (.A(tie_low_T13Y29), .B(tie_low_T13Y29), .X(2202));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9405  (.A(tie_low_T10Y26), .B(tie_low_T10Y26), .Y(2203));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9406  (.A(tie_low_T16Y24), .B(tie_low_T16Y24), .X(2204));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9407  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .X(2205));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9408  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .Y(2206));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9409  (.A(2203), .B(2206), .X(2207));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9410  (.A(tie_low_T12Y7), .B(tie_low_T12Y7), .X(2208));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9411  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(2209));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9412  (.A(tie_low_T7Y16), .B(tie_low_T7Y16), .Y(2210));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9413  (.A(tie_low_T7Y16), .B(tie_low_T7Y16), .X(2211));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9414  (.A(tie_low_T9Y16), .B(tie_low_T9Y16), .Y(2212));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9415  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(2213));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9416  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(2215));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9417  (.A(tie_low_T35Y60), .B(tie_low_T35Y60), .X(2216));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9418  (.A(tie_low_T15Y36), .B(tie_low_T15Y36), .Y(567));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9419  (.A(567), .Y(256));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9420  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .X(2217));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9421  (.A(2217), .Y(2218));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9422  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2219));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9423  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2220));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9424  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2221));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9425  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2222));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9426  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2223));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9427  (.A(286), .B(2203), .Y(2224));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9428  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(2225));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9429  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(2226));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9430  (.A(tie_low_T8Y18), .B(tie_low_T8Y18), .Y(2227));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9431  (.A(tie_low_T8Y16), .B(tie_low_T8Y16), .X(2228));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9432  (.A(2227), .B(2228), .Y(2229));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9433  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(2230));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9434  (.A(39), .B(2231), .X(2232));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9435  (.A(tie_low_T35Y70), .B(tie_low_T35Y70), .X(2233));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9436  (.A(tie_low_T15Y37), .B(tie_low_T15Y37), .Y(508));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9437  (.A(508), .Y(281));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9438  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .X(2234));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9439  (.A(2234), .Y(2235));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9440  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2236));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9441  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .X(2237));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9442  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2238));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9443  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .Y(2239));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9444  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2240));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9445  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .Y(2241));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9446  (.A(2241), .Y(2242));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9447  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .X(2243));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9448  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(2244));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9449  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(2245));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9450  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(2246));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9451  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .X(2247));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9452  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(2248));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9453  (.A(tie_low_T14Y16), .B(tie_low_T14Y16), .Y(2249));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9454  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(2251));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9455  (.A(tie_low_T35Y80), .B(tie_low_T35Y80), .X(2252));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9456  (.A(tie_low_T15Y41), .B(tie_low_T15Y41), .Y(1015));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9457  (.A(1015), .Y(305));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9458  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .X(2253));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9459  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(2254));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9460  (.A(2254), .Y(2255));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9461  (.A(tie_low_T13Y16), .B(tie_low_T13Y16), .Y(2256));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9462  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2257));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9463  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2258));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9464  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2259));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9465  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(2260));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9466  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .Y(2261));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9467  (.A(145), .B(2202), .X(2262));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9468  (.A(2261), .B(2262), .Y(2263));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9469  (.A(2263), .Y(2264));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9470  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(2265));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9471  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .X(2266));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9472  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(2267));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9473  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .X(2268));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9474  (.A(39), .B(2269), .X(2270));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9475  (.A(tie_low_T35Y89), .B(tie_low_T35Y89), .X(2271));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9476  (.A(tie_low_T15Y42), .B(tie_low_T15Y42), .Y(468));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9477  (.A(468), .Y(329));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9478  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .X(2272));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9479  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(2273));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9480  (.A(2273), .Y(2274));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9481  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(2275));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9482  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2276));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9483  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2277));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9484  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2278));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9485  (.A(tie_low_T14Y13), .B(tie_low_T14Y13), .X(2280));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9486  (.A(tie_low_T11Y27), .B(tie_low_T11Y27), .X(2281));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9487  (.A(tie_low_T10Y26), .B(tie_low_T10Y26), .Y(2282));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9488  (.A(tie_low_T12Y24), .B(tie_low_T12Y24), .X(2283));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9489  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .X(2284));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9490  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2285));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9491  (.A(2282), .B(2285), .X(2286));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9492  (.A(tie_low_T12Y7), .B(tie_low_T12Y7), .X(2287));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9493  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(2288));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9494  (.A(tie_low_T6Y16), .B(tie_low_T6Y16), .Y(2289));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9495  (.A(tie_low_T6Y16), .B(tie_low_T6Y16), .X(2290));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9496  (.A(tie_low_T8Y16), .B(tie_low_T8Y16), .Y(2291));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9497  (.A(tie_low_T14Y16), .B(tie_low_T14Y16), .Y(2292));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9498  (.A(tie_low_T0Y89), .B(tie_low_T0Y89), .Y(2293));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9499  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(2295));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9500  (.A(tie_low_T13Y34), .B(tie_low_T13Y34), .Y(352));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9501  (.A(tie_low_T14Y18), .B(tie_low_T14Y18), .X(2296));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9502  (.A(2296), .Y(2297));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9503  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2298));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9504  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2299));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9505  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2300));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9506  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2301));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9507  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2302));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9508  (.A(191), .B(2282), .Y(2303));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9509  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(2304));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9510  (.A(tie_low_T8Y22), .B(tie_low_T8Y22), .Y(2305));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9511  (.A(tie_low_T7Y17), .B(tie_low_T7Y17), .Y(2306));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9512  (.A(tie_low_T7Y16), .B(tie_low_T7Y16), .X(2307));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9513  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .Y(2308));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9514  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(2309));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9515  (.A(tie_low_T0Y51), .B(tie_low_T0Y51), .X(2311));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9516  (.A(tie_low_T3Y89), .B(tie_low_T3Y89), .X(2312));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9517  (.A(tie_low_T8Y41), .B(tie_low_T8Y41), .Y(1028));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9518  (.A(1028), .Y(375));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9519  (.A(tie_low_T14Y16), .B(tie_low_T14Y16), .X(2313));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9520  (.A(2313), .Y(2314));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9521  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2315));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9522  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .X(2316));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9523  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .X(2317));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9524  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2318));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9525  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2319));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9526  (.A(tie_low_T8Y21), .B(tie_low_T8Y21), .Y(2320));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9527  (.A(2320), .Y(2321));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9528  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(2322));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9529  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(2323));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9530  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(2324));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9531  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(2325));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9532  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .X(2326));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9533  (.A(2325), .B(2326), .Y(2327));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9534  (.A(tie_low_T14Y16), .B(tie_low_T14Y16), .Y(2328));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9535  (.A(39), .B(2329), .X(2330));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9536  (.A(tie_low_T7Y89), .B(tie_low_T7Y89), .X(2331));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9537  (.A(tie_low_T9Y39), .B(tie_low_T9Y39), .Y(1033));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9538  (.A(1033), .Y(398));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9539  (.A(tie_low_T14Y15), .B(tie_low_T14Y15), .X(2332));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9540  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(2333));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9541  (.A(2333), .Y(2334));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9542  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(2335));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9543  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .X(2336));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9544  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .Y(2337));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9545  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2338));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9546  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(2339));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9547  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .Y(2340));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9548  (.A(tie_low_T10Y27), .B(tie_low_T10Y27), .X(2341));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9549  (.A(tie_low_T10Y26), .B(tie_low_T10Y26), .Y(2342));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9550  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .X(2343));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9551  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(2344));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9552  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .Y(2345));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9553  (.A(tie_low_T14Y17), .B(tie_low_T14Y17), .Y(2346));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9554  (.A(tie_low_T21Y66), .B(tie_low_T21Y66), .Y(2348));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9555  (.A(tie_low_T11Y89), .B(tie_low_T11Y89), .Y(585));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9556  (.A(tie_low_T15Y45), .B(tie_low_T15Y45), .Y(419));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9557  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .X(2349));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9558  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(2350));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9559  (.A(2350), .Y(2351));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9560  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(2352));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9561  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2353));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9562  (.A(tie_low_T13Y14), .B(tie_low_T13Y14), .Y(2354));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9563  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2355));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9564  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .X(2356));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9565  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2357));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9566  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2358));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9567  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(2359));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9568  (.A(tie_low_T15Y6), .B(tie_low_T15Y6), .Y(2360));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9569  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2361));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9570  (.A(tie_low_T16Y6), .B(tie_low_T16Y6), .Y(2362));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9571  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2363));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9572  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2364));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9573  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(2365));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9574  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2366));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9575  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2367));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9576  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(2368));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9577  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2369));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9578  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2370));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9579  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(2371));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9580  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2372));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9581  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2373));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9582  (.A(tie_low_T15Y7), .B(tie_low_T15Y7), .Y(2374));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9583  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2375));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9584  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2376));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9585  (.A(tie_low_T15Y6), .B(tie_low_T15Y6), .Y(2377));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9586  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2378));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9587  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .X(2379));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9588  (.A(tie_low_T15Y6), .B(tie_low_T15Y6), .Y(2380));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9589  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .Y(482));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9590  (.A(tie_low_T7Y31), .B(tie_low_T7Y31), .X(2381));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9591  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2382));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9592  (.A(2220), .B(2381), .X(2383));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9593  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2384));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9594  (.A(2237), .B(2381), .X(2385));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9595  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2386));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9596  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2387));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9597  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2388));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9598  (.A(2256), .B(2381), .X(2389));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9599  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2390));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9600  (.A(2275), .B(2381), .X(2391));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9601  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2392));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9602  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2393));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9603  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2394));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9604  (.A(2299), .B(2381), .X(2395));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9605  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2396));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9606  (.A(2316), .B(2381), .X(2397));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9607  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2398));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9608  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2399));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9609  (.A(2335), .B(2381), .X(2400));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9610  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2401));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9611  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .Y(2402));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9612  (.A(2352), .B(2381), .X(2403));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9613  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2404));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9614  (.A(tie_low_T14Y11), .B(tie_low_T14Y11), .Y(2405));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9615  (.A(tie_low_T14Y10), .B(tie_low_T14Y10), .X(715));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9616  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .X(2406));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9617  (.A(2136), .B(2406), .Y(2407));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9618  (.A(2220), .B(2406), .X(2408));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9619  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2409));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9620  (.A(2237), .B(2406), .X(2410));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9621  (.A(714), .B(2406), .Y(2411));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9622  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2412));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9623  (.A(2256), .B(2406), .X(2413));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9624  (.A(746), .B(2406), .Y(2414));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9625  (.A(tie_low_T13Y13), .B(tie_low_T13Y13), .Y(2415));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9626  (.A(772), .B(2406), .Y(2416));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9627  (.A(2275), .B(2406), .X(2417));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9628  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2418));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9629  (.A(2299), .B(2406), .X(2419));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9630  (.A(804), .B(2406), .Y(2420));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9631  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2421));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9632  (.A(2316), .B(2406), .X(2422));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9633  (.A(833), .B(2406), .Y(2423));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9634  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2424));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9635  (.A(2335), .B(2406), .X(2425));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9636  (.A(862), .B(2406), .Y(2426));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9637  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2427));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9638  (.A(888), .B(2406), .Y(2428));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9639  (.A(2352), .B(2406), .X(2429));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9640  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2430));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9641  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .X(2431));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9642  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(2432));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9643  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(2433));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9644  (.A(tie_low_T13Y29), .B(tie_low_T13Y29), .Y(2434));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9645  (.A(tie_low_T13Y29), .B(tie_low_T13Y29), .X(2435));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9646  (.A(tie_low_T13Y29), .B(tie_low_T13Y29), .Y(2436));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9647  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(2437));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9648  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .X(2438));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9649  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(2439));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9650  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(2440));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9651  (.A(2440), .Y(2441));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9652  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(2442));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9653  (.A(tie_low_T11Y11), .B(tie_low_T11Y11), .Y(2443));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9654  (.A(2137), .B(2443), .Y(2444));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9655  (.A(2444), .Y(2445));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9656  (.A(tie_low_T13Y28), .B(tie_low_T13Y28), .Y(2446));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9657  (.A(2446), .Y(2447));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9658  (.A(tie_low_T10Y23), .B(tie_low_T10Y23), .Y(2448));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9659  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(2449));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9660  (.A(488), .B(2449), .X(469));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9661  (.A(469), .Y(542));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9662  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(2450));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9663  (.A(2450), .Y(466));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9664  (.A(2448), .B(466), .Y(2451));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9665  (.A(2447), .B(2451), .X(2452));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9666  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(2453));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9667  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(1113));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9668  (.A(1113), .Y(1517));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9669  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2454));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9670  (.A(472), .B(2454), .X(494));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9671  (.A(469), .B(494), .Y(2455));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9672  (.A(2455), .Y(501));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9673  (.A(tie_low_T9Y23), .B(tie_low_T9Y23), .X(476));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9674  (.A(tie_low_T14Y12), .B(tie_low_T14Y12), .X(2456));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9675  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .X(2457));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9676  (.A(472), .B(2457), .Y(2458));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9677  (.A(1254), .B(2458), .Y(2459));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9678  (.A(tie_low_T13Y17), .B(tie_low_T13Y17), .Y(2460));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9679  (.A(tie_low_T14Y14), .B(tie_low_T14Y14), .Y(2461));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9680  (.A(tie_low_T13Y15), .B(tie_low_T13Y15), .Y(2462));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9681  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2463));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9682  (.A(2463), .Y(2464));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9683  (.A(tie_low_T19Y66), .B(tie_low_T19Y66), .X(1404));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9684  (.A(1404), .Y(1387));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9685  (.A(tie_low_T13Y24), .B(tie_low_T13Y24), .Y(2465));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9686  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .X(2466));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9687  (.A(tie_low_T0Y30), .B(tie_low_T0Y30), .Y(2468));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9688  (.A(tie_low_T0Y30), .B(tie_low_T0Y30), .X(2092));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9689  (.A(tie_low_T8Y15), .B(tie_low_T8Y15), .X(2469));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9690  (.A(tie_low_T6Y22), .B(tie_low_T6Y22), .Y(2470));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9691  (.A(tie_low_T4Y16), .B(tie_low_T4Y16), .Y(2471));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9692  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .Y(2472));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9693  (.A(tie_low_T11Y13), .B(tie_low_T11Y13), .Y(2473));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9694  (.A(tie_low_T3Y19), .B(tie_low_T3Y19), .X(2474));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9695  (.A(2474), .Y(2475));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9696  (.A(tie_low_T15Y17), .B(tie_low_T15Y17), .X(2476));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9697  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .Y(2477));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9698  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(2478));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9699  (.A(2478), .Y(2479));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9700  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .Y(1455));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9701  (.A(1455), .Y(2480));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9702  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .X(2481));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9703  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .Y(2482));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9704  (.A(tie_low_T11Y13), .B(tie_low_T11Y13), .Y(2483));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9705  (.A(tie_low_T4Y18), .B(tie_low_T4Y18), .X(1349));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9706  (.A(1349), .Y(1174));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9707  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(2484));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9708  (.A(tie_low_T2Y20), .B(tie_low_T2Y20), .Y(1094));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9709  (.A(1094), .Y(1058));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9710  (.A(tie_low_T4Y27), .B(tie_low_T4Y27), .Y(450));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9711  (.A(450), .Y(1497));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9712  (.A(tie_low_T6Y23), .B(tie_low_T6Y23), .Y(1087));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9713  (.A(1087), .Y(1083));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9714  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .X(2485));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9715  (.A(tie_low_T15Y9), .B(tie_low_T15Y9), .Y(2486));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9716  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(2487));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9717  (.A(tie_low_T6Y26), .B(tie_low_T6Y26), .Y(1506));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9718  (.A(tie_low_T4Y28), .B(tie_low_T4Y28), .X(1049));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9719  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1046));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9720  (.A(tie_low_T2Y26), .B(tie_low_T2Y26), .Y(445));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9721  (.A(tie_low_T2Y37), .B(tie_low_T2Y37), .X(1040));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9722  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .X(2488));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9723  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .Y(2489));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9724  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(2490));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9725  (.A(2490), .Y(2491));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9726  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(2492));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9727  (.A(2492), .Y(2493));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9728  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .X(2494));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9729  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .Y(2495));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9730  (.A(tie_low_T11Y12), .B(tie_low_T11Y12), .Y(2496));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9731  (.A(tie_low_T3Y16), .B(tie_low_T3Y16), .X(2497));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9732  (.A(2497), .Y(1097));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9733  (.A(tie_low_T3Y21), .B(tie_low_T3Y21), .Y(2498));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9734  (.A(tie_low_T5Y27), .B(tie_low_T5Y27), .X(1055));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9735  (.A(1055), .Y(1431));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9736  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .X(2499));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9737  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .Y(2500));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9738  (.A(tie_low_T11Y13), .B(tie_low_T11Y13), .Y(2501));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9739  (.A(tie_low_T4Y19), .B(tie_low_T4Y19), .X(2502));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9740  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .X(2503));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9741  (.A(tie_low_T15Y10), .B(tie_low_T15Y10), .Y(2504));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9742  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(2505));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9743  (.A(2505), .Y(2506));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9744  (.A(tie_low_T6Y25), .B(tie_low_T6Y25), .Y(1061));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9745  (.A(tie_low_T3Y23), .B(tie_low_T3Y23), .Y(1069));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9746  (.A(tie_low_T4Y25), .B(tie_low_T4Y25), .X(1395));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9747  (.A(tie_low_T7Y28), .B(tie_low_T7Y28), .X(1047));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9748  (.A(tie_low_T15Y30), .B(tie_low_T15Y30), .X(2507));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9749  (.A(tie_low_T6Y32), .B(tie_low_T6Y32), .X(2508));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9750  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(2509));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9751  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2510));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9752  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(1076));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9753  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .X(1101));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9754  (.A(tie_low_T8Y31), .B(tie_low_T8Y31), .X(2511));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9755  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(2512));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9756  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(2513));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9757  (.A(tie_low_T6Y24), .B(tie_low_T6Y24), .Y(1460));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9758  (.A(tie_low_T4Y28), .B(tie_low_T4Y28), .Y(440));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9759  (.A(440), .Y(2514));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9760  (.A(tie_low_T5Y34), .B(tie_low_T5Y34), .X(1412));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9761  (.A(tie_low_T7Y32), .B(tie_low_T7Y32), .X(2515));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9762  (.A(tie_low_T6Y30), .B(tie_low_T6Y30), .X(2516));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9763  (.A(2513), .B(2516), .Y(2517));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9764  (.A(tie_low_T17Y31), .B(tie_low_T17Y31), .Y(2518));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9765  (.A(tie_low_T5Y34), .B(tie_low_T5Y34), .Y(2519));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9766  (.A(tie_low_T7Y32), .B(tie_low_T7Y32), .X(2520));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9767  (.A(tie_low_T6Y30), .B(tie_low_T6Y30), .X(2521));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9768  (.A(tie_low_T14Y20), .B(tie_low_T14Y20), .Y(2522));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9769  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2523));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9770  (.A(tie_low_T4Y37), .B(tie_low_T4Y37), .Y(1477));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9771  (.A(tie_low_T5Y32), .B(tie_low_T5Y32), .X(2524));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9772  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(2525));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9773  (.A(tie_low_T17Y31), .B(tie_low_T17Y31), .Y(2526));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9774  (.A(tie_low_T5Y32), .B(tie_low_T5Y32), .X(2527));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9775  (.A(tie_low_T13Y21), .B(tie_low_T13Y21), .Y(2528));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9776  (.A(tie_low_T13Y24), .B(tie_low_T13Y24), .Y(2529));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9777  (.A(tie_low_T5Y35), .B(tie_low_T5Y35), .X(1050));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9778  (.A(tie_low_T6Y32), .B(tie_low_T6Y32), .X(2530));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9779  (.A(tie_low_T12Y19), .B(tie_low_T12Y19), .Y(2531));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9780  (.A(tie_low_T18Y32), .B(tie_low_T18Y32), .Y(2532));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9781  (.A(tie_low_T6Y32), .B(tie_low_T6Y32), .X(2533));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9782  (.A(tie_low_T14Y22), .B(tie_low_T14Y22), .Y(2534));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9783  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2535));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9784  (.A(tie_low_T3Y35), .B(tie_low_T3Y35), .X(1413));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9785  (.A(1413), .Y(2536));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9786  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(2537));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9787  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(2538));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9788  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2539));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9789  (.A(tie_low_T4Y27), .B(tie_low_T4Y27), .X(2540));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9790  (.A(tie_low_T4Y27), .B(tie_low_T4Y27), .X(2541));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9791  (.A(tie_low_T6Y31), .B(tie_low_T6Y31), .X(1463));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9792  (.A(tie_low_T15Y30), .B(tie_low_T15Y30), .X(2542));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9793  (.A(tie_low_T16Y20), .B(tie_low_T16Y20), .Y(2543));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9794  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2544));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9795  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1072));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9796  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(1085));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9797  (.A(tie_low_T4Y29), .B(tie_low_T4Y29), .X(2545));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9798  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .Y(2546));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9799  (.A(tie_low_T14Y33), .B(tie_low_T14Y33), .X(2547));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9800  (.A(2547), .Y(2548));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9801  (.A(tie_low_T7Y29), .B(tie_low_T7Y29), .Y(2549));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9802  (.A(tie_low_T5Y35), .B(tie_low_T5Y35), .X(2550));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9803  (.A(tie_low_T5Y36), .B(tie_low_T5Y36), .X(2551));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9804  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(2552));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9805  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .X(1464));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9806  (.A(tie_low_T15Y31), .B(tie_low_T15Y31), .X(2553));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9807  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2554));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9808  (.A(tie_low_T16Y20), .B(tie_low_T16Y20), .Y(2555));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9809  (.A(tie_low_T3Y23), .B(tie_low_T3Y23), .Y(1062));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9810  (.A(1062), .Y(2556));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9811  (.A(tie_low_T4Y28), .B(tie_low_T4Y28), .X(1052));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9812  (.A(1052), .Y(1043));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9813  (.A(tie_low_T4Y29), .B(tie_low_T4Y29), .X(1041));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9814  (.A(tie_low_T5Y27), .B(tie_low_T5Y27), .X(2557));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9815  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(2558));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9816  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .X(1393));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9817  (.A(tie_low_T4Y24), .B(tie_low_T4Y24), .X(2559));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9818  (.A(tie_low_T5Y27), .B(tie_low_T5Y27), .X(2560));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9819  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(1484));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9820  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(1073));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9821  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(1088));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9822  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .X(1495));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9823  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .X(2561));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9824  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(2562));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9825  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(2563));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9826  (.A(tie_low_T15Y30), .B(tie_low_T15Y30), .Y(2564));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9827  (.A(tie_low_T12Y27), .B(tie_low_T12Y27), .Y(2565));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9828  (.A(2565), .Y(2566));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9829  (.A(tie_low_T15Y28), .B(tie_low_T15Y28), .Y(2567));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9830  (.A(tie_low_T13Y21), .B(tie_low_T13Y21), .Y(2568));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9831  (.A(tie_low_T8Y27), .B(tie_low_T8Y27), .Y(2569));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9832  (.A(39), .B(2569), .Y(2570));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9833  (.A(tie_low_T12Y18), .B(tie_low_T12Y18), .Y(2571));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9834  (.A(tie_low_T4Y37), .B(tie_low_T4Y37), .Y(1456));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9835  (.A(tie_low_T7Y28), .B(tie_low_T7Y28), .X(2572));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9836  (.A(tie_low_T5Y32), .B(tie_low_T5Y32), .X(2573));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9837  (.A(2571), .B(2573), .Y(2574));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9838  (.A(1886), .B(2570), .Y(2575));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9839  (.A(tie_low_T14Y9), .B(tie_low_T14Y9), .Y(2576));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9840  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(2577));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9841  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2578));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9842  (.A(tie_low_T5Y32), .B(tie_low_T5Y32), .X(1473));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9843  (.A(tie_low_T5Y35), .B(tie_low_T5Y35), .X(2579));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9844  (.A(tie_low_T9Y30), .B(tie_low_T9Y30), .X(2580));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9845  (.A(tie_low_T9Y28), .B(tie_low_T9Y28), .Y(2581));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9846  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(2582));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9847  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2583));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9848  (.A(tie_low_T15Y17), .B(tie_low_T15Y17), .Y(2584));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9849  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .X(1397));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9850  (.A(tie_low_T15Y30), .B(tie_low_T15Y30), .X(2585));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9851  (.A(tie_low_T12Y22), .B(tie_low_T12Y22), .Y(2586));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9852  (.A(tie_low_T15Y18), .B(tie_low_T15Y18), .Y(2587));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9853  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2588));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9854  (.A(tie_low_T7Y30), .B(tie_low_T7Y30), .Y(2589));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9855  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(2590));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9856  (.A(tie_low_T12Y20), .B(tie_low_T12Y20), .Y(2591));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9857  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .Y(2592));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9858  (.A(tie_low_T15Y29), .B(tie_low_T15Y29), .Y(2593));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9859  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .Y(2594));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9860  (.A(tie_low_T13Y33), .B(tie_low_T13Y33), .X(2595));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9861  (.A(tie_low_T12Y26), .B(tie_low_T12Y26), .X(2596));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9862  (.A(tie_low_T16Y15), .B(tie_low_T16Y15), .Y(2597));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9863  (.A(tie_low_T4Y27), .B(tie_low_T4Y27), .Y(1056));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9864  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(1064));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9865  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1219));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9866  (.A(tie_low_T7Y27), .B(tie_low_T7Y27), .X(1095));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9867  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(2598));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9868  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(2599));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9869  (.A(2599), .Y(1438));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9870  (.A(tie_low_T4Y26), .B(tie_low_T4Y26), .X(2600));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9871  (.A(tie_low_T4Y30), .B(tie_low_T4Y30), .X(2601));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9872  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(2602));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9873  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(2603));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9874  (.A(tie_low_T13Y19), .B(tie_low_T13Y19), .X(2604));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9875  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .Y(2605));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9876  (.A(2605), .Y(2606));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9877  (.A(tie_low_T13Y19), .B(tie_low_T13Y19), .X(2607));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9878  (.A(tie_low_T8Y30), .B(tie_low_T8Y30), .Y(2608));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9879  (.A(tie_low_T6Y29), .B(tie_low_T6Y29), .Y(2609));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9880  (.A(2609), .Y(2610));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9881  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(2611));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9882  (.A(tie_low_T6Y25), .B(tie_low_T6Y25), .X(1445));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9883  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(2612));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9884  (.A(tie_low_T5Y36), .B(tie_low_T5Y36), .X(1436));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9885  (.A(tie_low_T4Y28), .B(tie_low_T4Y28), .X(2613));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9886  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .Y(2614));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9887  (.A(2614), .Y(2615));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9888  (.A(tie_low_T4Y27), .B(tie_low_T4Y27), .X(1389));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9889  (.A(tie_low_T5Y28), .B(tie_low_T5Y28), .X(1428));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9890  (.A(tie_low_T5Y31), .B(tie_low_T5Y31), .X(1479));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9891  (.A(1479), .Y(1406));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9892  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(2616));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9893  (.A(tie_low_T5Y29), .B(tie_low_T5Y29), .Y(2617));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9894  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(2618));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9895  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .X(2619));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9896  (.A(tie_low_T4Y26), .B(tie_low_T4Y26), .X(2620));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9897  (.A(tie_low_T5Y27), .B(tie_low_T5Y27), .Y(2621));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9898  (.A(2621), .Y(2622));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9899  (.A(tie_low_T5Y30), .B(tie_low_T5Y30), .Y(2623));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9900  (.A(tie_low_T6Y28), .B(tie_low_T6Y28), .X(2624));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9901  (.A(tie_low_T12Y21), .B(tie_low_T12Y21), .Y(2625));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9902  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(2626));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9903  (.A(tie_low_T11Y22), .B(tie_low_T11Y22), .X(2627));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9904  (.A(tie_low_T13Y19), .B(tie_low_T13Y19), .Y(2628));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9905  (.A(2628), .Y(2629));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9906  (.A(tie_low_T7Y20), .B(tie_low_T7Y20), .X(2630));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9907  (.A(tie_low_T10Y17), .B(tie_low_T10Y17), .X(621));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9908  (.A(tie_low_T6Y17), .B(tie_low_T6Y17), .X(172));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9909  (.A(172), .Y(148));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9910  (.A(tie_low_T14Y29), .B(tie_low_T14Y29), .X(2631));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9911  (.A(tie_low_T14Y29), .B(tie_low_T14Y29), .Y(2632));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9912  (.A(tie_low_T11Y24), .B(tie_low_T11Y24), .Y(1184));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9913  (.A(tie_low_T10Y22), .B(tie_low_T10Y22), .Y(1331));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9914  (.A(tie_low_T9Y22), .B(tie_low_T9Y22), .Y(2633));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9915  (.A(tie_low_T9Y15), .B(tie_low_T9Y15), .Y(2634));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9916  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(264));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9917  (.A(264), .Y(287));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9918  (.A(488), .B(2453), .X(2635));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9919  (.A(tie_low_T8Y21), .B(tie_low_T8Y21), .Y(2636));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9920  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .X(2637));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9921  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .X(2638));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9922  (.A(tie_low_T0Y0), .B(tie_low_T0Y0), .Y(1578));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9923  (.A(tie_low_T8Y15), .B(tie_low_T8Y15), .X(2639));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9924  (.A(2639), .Y(2640));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9925  (.A(tie_low_T12Y16), .B(tie_low_T12Y16), .X(2641));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9926  (.A(2153), .B(609), .X(631));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9927  (.A(488), .B(631), .X(2642));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9928  (.A(2641), .B(2642), .Y(1115));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9929  (.A(614), .B(631), .X(1126));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9930  (.A(1126), .Y(2643));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9931  (.A(tie_low_T11Y21), .B(tie_low_T11Y21), .X(650));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9932  (.A(tie_low_T8Y17), .B(tie_low_T8Y17), .X(1295));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9933  (.A(1295), .Y(1262));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9934  (.A(666), .B(615), .Y(691));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9935  (.A(tie_low_T9Y20), .B(tie_low_T9Y20), .Y(1201));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9936  (.A(tie_low_T9Y18), .B(tie_low_T9Y18), .Y(1144));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9937  (.A(650), .B(1144), .X(2644));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9938  (.A(tie_low_T7Y28), .B(tie_low_T7Y28), .X(2645));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9939  (.A(tie_low_T4Y37), .B(tie_low_T4Y37), .X(2646));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9940  (.A(614), .B(2453), .X(2647));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9941  (.A(tie_low_T10Y20), .B(tie_low_T10Y20), .Y(1119));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9942  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .X(146));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9943  (.A(tie_low_T9Y17), .B(tie_low_T9Y17), .X(150));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9944  (.A(150), .Y(199));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9945  (.A(tie_low_T7Y21), .B(tie_low_T7Y21), .Y(2648));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9946  (.A(tie_low_T9Y21), .B(tie_low_T9Y21), .X(1141));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9947  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(2649));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9948  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .X(2650));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9949  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(254));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9950  (.A(tie_low_T9Y25), .B(tie_low_T9Y25), .X(143));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9951  (.A(tie_low_T10Y25), .B(tie_low_T10Y25), .Y(2651));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9952  (.A(516), .B(146), .Y(2652));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9953  (.A(tie_low_T9Y24), .B(tie_low_T9Y24), .X(2653));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9954  (.A(2653), .Y(153));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9955  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(2654));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9956  (.A(tie_low_T7Y17), .B(tie_low_T7Y17), .X(681));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9957  (.A(tie_low_T10Y15), .B(tie_low_T10Y15), .Y(2655));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9958  (.A(2655), .Y(2656));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9959  (.A(2652), .B(2656), .Y(2657));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9960  (.A(2657), .Y(2658));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9961  (.A(tie_low_T5Y36), .B(tie_low_T5Y36), .Y(2659));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9962  (.A(tie_low_T0Y47), .B(tie_low_T0Y47), .Y(2660));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9963  (.A(2660), .Y(2661));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9964  (.A(tie_low_T2Y43), .B(tie_low_T2Y43), .X(2662));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9965  (.A(tie_low_T0Y47), .B(tie_low_T0Y47), .Y(2663));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9966  (.A(39), .B(2663), .Y(2664));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9967  (.A(675), .B(39), .X(2665));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9968  (.A(2664), .B(2665), .Y(2666));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9969  (.A(2666), .Y(2667));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9970  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(2668));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9971  (.A(286), .B(146), .Y(2669));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9972  (.A(tie_low_T15Y11), .B(tie_low_T15Y11), .Y(2670));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9973  (.A(286), .B(148), .Y(2671));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9974  (.A(2671), .Y(729));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9975  (.A(tie_low_T12Y13), .B(tie_low_T12Y13), .Y(2673));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9976  (.A(tie_low_T13Y12), .B(tie_low_T13Y12), .Y(2674));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9977  (.A(2669), .B(2671), .Y(2675));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9978  (.A(2674), .B(2675), .X(2676));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9979  (.A(2676), .Y(2677));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9980  (.A(tie_low_T5Y37), .B(tie_low_T5Y37), .Y(2678));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9981  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(2679));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9982  (.A(2679), .Y(132));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9983  (.A(tie_low_T2Y44), .B(tie_low_T2Y44), .X(2680));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9984  (.A(tie_low_T0Y48), .B(tie_low_T0Y48), .Y(2681));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9985  (.A(39), .B(2681), .Y(2682));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9986  (.A(39), .B(721), .X(2683));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9987  (.A(2682), .B(2683), .Y(2684));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9988  (.A(2684), .Y(2685));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9989  (.A(tie_low_T11Y25), .B(tie_low_T11Y25), .Y(130));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9990  (.A(518), .B(146), .Y(2686));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9991  (.A(2686), .Y(127));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9992  (.A(tie_low_T15Y12), .B(tie_low_T15Y12), .Y(2687));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9993  (.A(tie_low_T6Y17), .B(tie_low_T6Y17), .X(2688));
  sky130_fd_sc_hd__clkinv_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9994  (.A(2688), .Y(124));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9995  (.A(tie_low_T19Y29), .B(tie_low_T19Y29), .Y(2689));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9996  (.A(tie_low_T16Y12), .B(tie_low_T16Y12), .X(2691));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9997  (.A(tie_low_T15Y20), .B(tie_low_T15Y20), .Y(2692));
  sky130_fd_sc_hd__or2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9998  (.A(tie_low_T10Y19), .B(tie_low_T10Y19), .X(2693));
  sky130_fd_sc_hd__nand2_2 \$abc$9276$auto$blifparse.cc:396:parse_blif$9999  (.A(tie_low_T12Y15), .B(tie_low_T12Y15), .Y(125));
  sky130_fd_sc_hd__conb_1 \$auto$hilomap.cc:40:hilomap_worker$12031  (.HI(2694));
  sky130_fd_sc_hd__conb_1 \$auto$hilomap.cc:40:hilomap_worker$8815  (.HI(60));
  sky130_fd_sc_hd__conb_1 \$auto$hilomap.cc:48:hilomap_worker$8817  (.LO(44));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11708  (.A(531), .Y(2695));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11709  (.A(577), .Y(2696));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11710  (.A(2110), .Y(2697));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11711  (.A(2121), .Y(2698));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11712  (.A(44), .Y(2699));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11713  (.A(60), .Y(2700));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11714  (.A(60), .Y(2701));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11715  (.A(44), .Y(2702));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11716  (.A(60), .Y(2703));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11717  (.A(44), .Y(2704));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11718  (.A(60), .Y(2705));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11719  (.A(60), .Y(2706));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11720  (.A(44), .Y(2707));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11721  (.A(60), .Y(2708));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11722  (.A(44), .Y(2709));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11723  (.A(44), .Y(2710));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11724  (.A(44), .Y(2711));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11725  (.A(60), .Y(2712));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11726  (.A(44), .Y(2713));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11727  (.A(60), .Y(2714));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11728  (.A(44), .Y(2715));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11729  (.A(44), .Y(2716));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11730  (.A(60), .Y(2717));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11731  (.A(44), .Y(2718));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11732  (.A(44), .Y(2719));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11733  (.A(60), .Y(2720));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11734  (.A(44), .Y(2721));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11735  (.A(44), .Y(2722));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11736  (.A(60), .Y(2723));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11737  (.A(44), .Y(2724));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11738  (.A(44), .Y(2725));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11739  (.A(60), .Y(2726));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11740  (.A(60), .Y(2727));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11741  (.A(44), .Y(2728));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11742  (.A(44), .Y(2729));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11743  (.A(44), .Y(2730));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11744  (.A(60), .Y(2731));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11745  (.A(60), .Y(2732));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11746  (.A(44), .Y(2733));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11747  (.A(44), .Y(2734));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11748  (.A(60), .Y(2735));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11749  (.A(60), .Y(2736));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11750  (.A(60), .Y(2737));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11751  (.A(44), .Y(2738));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11752  (.A(60), .Y(2739));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11753  (.A(44), .Y(2740));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11754  (.A(2741), .Y(2742));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11755  (.A(60), .Y(2743));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11756  (.A(44), .Y(2744));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11757  (.A(44), .Y(2745));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11758  (.A(44), .Y(2746));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11759  (.A(60), .Y(2747));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11760  (.A(44), .Y(2748));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11761  (.A(44), .Y(2749));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11762  (.A(60), .Y(2750));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11763  (.A(44), .Y(2751));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11764  (.A(60), .Y(2752));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11765  (.A(60), .Y(2753));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11766  (.A(44), .Y(2754));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11767  (.A(44), .Y(2755));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11768  (.A(60), .Y(2756));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11769  (.A(44), .Y(2757));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11770  (.A(60), .Y(2758));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11771  (.A(60), .Y(2759));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11772  (.A(44), .Y(2760));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11773  (.A(60), .Y(2761));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11774  (.A(44), .Y(2762));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11775  (.A(44), .Y(2763));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11776  (.A(60), .Y(2764));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11777  (.A(60), .Y(2765));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11778  (.A(44), .Y(2766));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11779  (.A(60), .Y(2767));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11780  (.A(60), .Y(2768));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11781  (.A(60), .Y(2769));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11782  (.A(44), .Y(2770));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11783  (.A(60), .Y(2771));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11784  (.A(44), .Y(2772));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11785  (.A(60), .Y(2773));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11786  (.A(60), .Y(2774));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11787  (.A(44), .Y(2775));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11788  (.A(44), .Y(2776));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11789  (.A(60), .Y(2777));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11790  (.A(44), .Y(2778));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11791  (.A(60), .Y(2779));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11792  (.A(44), .Y(2780));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11793  (.A(44), .Y(2781));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11794  (.A(44), .Y(2782));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11795  (.A(60), .Y(2783));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11796  (.A(44), .Y(2784));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11797  (.A(60), .Y(2785));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11798  (.A(60), .Y(2786));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11799  (.A(60), .Y(2787));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11800  (.A(60), .Y(2788));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11801  (.A(44), .Y(2789));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11802  (.A(44), .Y(2790));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11803  (.A(60), .Y(2791));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11804  (.A(44), .Y(2792));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11805  (.A(60), .Y(2793));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11806  (.A(60), .Y(2794));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11807  (.A(44), .Y(2795));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11808  (.A(44), .Y(2796));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11809  (.A(60), .Y(2797));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11810  (.A(60), .Y(2798));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11811  (.A(44), .Y(2799));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11812  (.A(60), .Y(2800));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11813  (.A(60), .Y(2801));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11814  (.A(60), .Y(2802));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11815  (.A(44), .Y(2803));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11816  (.A(44), .Y(2804));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11817  (.A(44), .Y(2805));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11818  (.A(60), .Y(2806));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11819  (.A(60), .Y(2807));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11820  (.A(60), .Y(2808));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11821  (.A(44), .Y(2809));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11822  (.A(60), .Y(2810));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11823  (.A(60), .Y(2811));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11824  (.A(44), .Y(2812));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11825  (.A(60), .Y(2813));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11826  (.A(60), .Y(2814));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11827  (.A(44), .Y(2815));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11828  (.A(44), .Y(2816));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11829  (.A(44), .Y(2817));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11830  (.A(44), .Y(2818));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11831  (.A(44), .Y(2819));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11832  (.A(44), .Y(2820));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11833  (.A(60), .Y(2821));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11834  (.A(60), .Y(2822));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11835  (.A(60), .Y(2823));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11836  (.A(60), .Y(2824));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11837  (.A(60), .Y(2825));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11838  (.A(60), .Y(2826));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11839  (.A(44), .Y(2827));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11840  (.A(44), .Y(2828));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11841  (.A(60), .Y(2829));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11842  (.A(44), .Y(2830));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11843  (.A(44), .Y(2831));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11844  (.A(44), .Y(2832));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11845  (.A(60), .Y(2833));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11846  (.A(44), .Y(2834));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11847  (.A(60), .Y(2835));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11848  (.A(60), .Y(2836));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11849  (.A(60), .Y(2837));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11850  (.A(44), .Y(2838));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11851  (.A(60), .Y(2839));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11852  (.A(60), .Y(2840));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11853  (.A(44), .Y(2841));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11854  (.A(60), .Y(2842));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11855  (.A(44), .Y(2843));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11856  (.A(44), .Y(2844));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11857  (.A(44), .Y(2845));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11858  (.A(60), .Y(2846));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11859  (.A(44), .Y(2847));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11860  (.A(60), .Y(2848));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11861  (.A(44), .Y(2849));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11862  (.A(60), .Y(2850));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11863  (.A(60), .Y(2851));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11864  (.A(44), .Y(2852));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11865  (.A(44), .Y(2853));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11866  (.A(60), .Y(2854));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11867  (.A(44), .Y(2855));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11868  (.A(60), .Y(2856));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11869  (.A(44), .Y(2857));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11870  (.A(44), .Y(2858));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11871  (.A(44), .Y(2859));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11872  (.A(60), .Y(2860));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11873  (.A(44), .Y(2861));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11874  (.A(44), .Y(2862));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11875  (.A(44), .Y(2863));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11876  (.A(44), .Y(2864));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11877  (.A(44), .Y(2865));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11878  (.A(60), .Y(2866));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11879  (.A(44), .Y(2867));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11880  (.A(60), .Y(2868));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11881  (.A(60), .Y(2869));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11882  (.A(60), .Y(2870));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11883  (.A(60), .Y(2871));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11884  (.A(44), .Y(2872));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11885  (.A(44), .Y(2873));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11886  (.A(60), .Y(2874));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11887  (.A(1196), .Y(2875));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11888  (.A(562), .Y(2876));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11889  (.A(44), .Y(2877));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11890  (.A(1196), .Y(2878));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11891  (.A(2879), .Y(2880));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11892  (.A(44), .Y(2881));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11893  (.A(60), .Y(2882));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11894  (.A(44), .Y(2883));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11895  (.A(44), .Y(2884));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11896  (.A(60), .Y(2885));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11897  (.A(60), .Y(2886));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11898  (.A(44), .Y(2887));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11899  (.A(44), .Y(2888));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11900  (.A(44), .Y(2889));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11901  (.A(44), .Y(2890));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11902  (.A(60), .Y(2891));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11903  (.A(44), .Y(2892));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11904  (.A(44), .Y(2893));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11905  (.A(44), .Y(2894));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11906  (.A(44), .Y(2895));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11907  (.A(44), .Y(2896));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11908  (.A(60), .Y(2897));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11909  (.A(44), .Y(2898));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11910  (.A(44), .Y(2899));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11911  (.A(44), .Y(2900));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11912  (.A(60), .Y(2901));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11913  (.A(60), .Y(2902));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11914  (.A(44), .Y(2903));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11915  (.A(60), .Y(2904));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11916  (.A(60), .Y(2905));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11917  (.A(60), .Y(2906));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11918  (.A(60), .Y(2907));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11919  (.A(60), .Y(2908));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11920  (.A(60), .Y(2909));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11921  (.A(60), .Y(2910));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11922  (.A(60), .Y(2911));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11923  (.A(60), .Y(2912));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11924  (.A(60), .Y(2913));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11925  (.A(60), .Y(2914));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11926  (.A(60), .Y(2915));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11927  (.A(60), .Y(2916));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11928  (.A(675), .Y(2917));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11929  (.A(721), .Y(2918));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11930  (.A(138), .Y(2919));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11931  (.A(142), .Y(2920));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11932  (.A(167), .Y(2921));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11933  (.A(189), .Y(2922));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11934  (.A(211), .Y(2923));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11935  (.A(232), .Y(2924));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11936  (.A(516), .Y(2925));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11937  (.A(286), .Y(2926));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11938  (.A(518), .Y(2927));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11939  (.A(145), .Y(2928));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11940  (.A(169), .Y(2929));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11941  (.A(191), .Y(2930));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11942  (.A(213), .Y(2931));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11943  (.A(234), .Y(2932));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11944  (.A(516), .Y(2933));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11945  (.A(286), .Y(2934));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11946  (.A(518), .Y(2935));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11947  (.A(145), .Y(2936));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11948  (.A(169), .Y(2937));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11949  (.A(191), .Y(2938));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11950  (.A(213), .Y(2939));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11951  (.A(234), .Y(2940));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11952  (.A(258), .Y(2941));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11953  (.A(283), .Y(2942));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11954  (.A(307), .Y(2943));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11955  (.A(331), .Y(2944));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11956  (.A(355), .Y(2945));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11957  (.A(378), .Y(2946));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11958  (.A(400), .Y(2947));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11959  (.A(421), .Y(2948));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11960  (.A(516), .Y(2949));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11961  (.A(286), .Y(2950));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11962  (.A(518), .Y(2951));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11963  (.A(145), .Y(2952));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11964  (.A(169), .Y(2953));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11965  (.A(191), .Y(2954));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11966  (.A(213), .Y(2955));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11967  (.A(234), .Y(2956));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11968  (.A(256), .Y(2957));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11969  (.A(281), .Y(2958));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11970  (.A(305), .Y(2959));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11971  (.A(329), .Y(2960));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11972  (.A(352), .Y(2961));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11973  (.A(375), .Y(2962));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11974  (.A(398), .Y(2963));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11975  (.A(419), .Y(2964));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11976  (.A(234), .Y(2965));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11977  (.A(44), .Y(45));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11978  (.A(44), .Y(54));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11979  (.A(44), .Y(55));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11980  (.A(44), .Y(56));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11981  (.A(44), .Y(57));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11982  (.A(44), .Y(58));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11983  (.A(44), .Y(59));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11984  (.A(60), .Y(61));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11985  (.A(60), .Y(62));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11986  (.A(60), .Y(63));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11987  (.A(44), .Y(46));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11988  (.A(60), .Y(64));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11989  (.A(60), .Y(65));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11990  (.A(60), .Y(66));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11991  (.A(60), .Y(67));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11992  (.A(44), .Y(68));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11993  (.A(44), .Y(69));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11994  (.A(44), .Y(70));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11995  (.A(44), .Y(71));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11996  (.A(44), .Y(72));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11997  (.A(44), .Y(73));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11998  (.A(44), .Y(47));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$11999  (.A(44), .Y(74));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12000  (.A(44), .Y(75));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12001  (.A(44), .Y(76));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12002  (.A(60), .Y(77));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12003  (.A(60), .Y(78));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12004  (.A(60), .Y(79));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12005  (.A(60), .Y(80));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12006  (.A(60), .Y(81));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12007  (.A(60), .Y(82));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12008  (.A(60), .Y(83));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12009  (.A(44), .Y(48));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12010  (.A(44), .Y(49));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12011  (.A(44), .Y(50));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12012  (.A(44), .Y(51));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12013  (.A(44), .Y(52));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12014  (.A(44), .Y(53));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12015  (.A(44), .Y(100));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12016  (.A(44), .Y(101));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12017  (.A(44), .Y(102));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12018  (.A(44), .Y(103));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12019  (.A(44), .Y(104));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12020  (.A(44), .Y(105));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12021  (.A(44), .Y(106));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12022  (.A(44), .Y(107));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12023  (.A(44), .Y(117));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12024  (.A(44), .Y(118));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12025  (.A(44), .Y(119));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12026  (.A(44), .Y(120));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12027  (.A(44), .Y(121));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12028  (.A(44), .Y(122));
  sky130_fd_sc_hd__clkbuf_4 \$auto$insbuf.cc:97:execute$12029  (.A(44), .Y(123));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4105  (.CLK(clk_cts_n6), .D(2223), .Q(597), .Q_N(2966), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4106  (.CLK(clk_cts_n6), .D(2240), .Q(2134), .Q_N(2967), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4107  (.CLK(clk_cts_n4), .D(2259), .Q(739), .Q_N(2968), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4108  (.CLK(clk_cts_n4), .D(2278), .Q(768), .Q_N(2969), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4109  (.CLK(clk_cts_n4), .D(2302), .Q(797), .Q_N(2970), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4110  (.CLK(clk_cts_n4), .D(2319), .Q(826), .Q_N(2971), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4111  (.CLK(clk_cts_n6), .D(2338), .Q(855), .Q_N(2972), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4112  (.CLK(clk_cts_n0), .D(2355), .Q(884), .Q_N(2973), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4907  (.CLK(clk_cts_n4), .D(2359), .Q(2135), .Q_N(2974), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4908  (.CLK(clk_cts_n0), .D(2362), .Q(707), .Q_N(2975), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4909  (.CLK(clk_cts_n0), .D(2365), .Q(736), .Q_N(2976), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4910  (.CLK(clk_cts_n0), .D(2368), .Q(766), .Q_N(2977), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4911  (.CLK(clk_cts_n0), .D(2371), .Q(795), .Q_N(2978), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4912  (.CLK(clk_cts_n0), .D(2374), .Q(824), .Q_N(2979), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4913  (.CLK(clk_cts_n4), .D(2377), .Q(853), .Q_N(2980), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4914  (.CLK(clk_cts_n6), .D(2380), .Q(882), .Q_N(2981), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4931  (.CLK(clk_cts_n0), .D(2384), .Q(590), .Q_N(2982), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4932  (.CLK(clk_cts_n4), .D(2387), .Q(711), .Q_N(2983), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4933  (.CLK(clk_cts_n0), .D(2390), .Q(743), .Q_N(2984), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4934  (.CLK(clk_cts_n4), .D(2393), .Q(775), .Q_N(2985), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4935  (.CLK(clk_cts_n0), .D(2396), .Q(801), .Q_N(2986), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4936  (.CLK(clk_cts_n0), .D(2399), .Q(830), .Q_N(2987), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4937  (.CLK(clk_cts_n0), .D(2402), .Q(859), .Q_N(2988), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4938  (.CLK(clk_cts_n0), .D(2405), .Q(891), .Q_N(2989), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4979  (.CLK(clk_cts_n0), .D(2409), .Q(2136), .Q_N(2990), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4980  (.CLK(clk_cts_n0), .D(2412), .Q(714), .Q_N(2991), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4981  (.CLK(clk_cts_n0), .D(2415), .Q(746), .Q_N(2992), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4982  (.CLK(clk_cts_n4), .D(2418), .Q(772), .Q_N(2993), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4983  (.CLK(clk_cts_n6), .D(2421), .Q(804), .Q_N(2994), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4984  (.CLK(clk_cts_n0), .D(2424), .Q(833), .Q_N(2995), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4985  (.CLK(clk_cts_n4), .D(2427), .Q(862), .Q_N(2996), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$4986  (.CLK(clk_cts_n0), .D(2430), .Q(888), .Q_N(2997), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5134  (.CLK(clk_cts_n4), .D(2464), .Q(2110), .Q_N(1251), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5135  (.CLK(clk_cts_n0), .D(1992), .Q(1988), .Q_N(2690), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5136  (.CLK(clk_cts_n1), .D(38), .Q(2998), .Q_N(1985), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5137  (.CLK(clk_cts_n2), .D(2509), .Q(462), .Q_N(2181), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5138  (.CLK(clk_cts_n0), .D(2512), .Q(2043), .Q_N(2999), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5139  (.CLK(clk_cts_n0), .D(2517), .Q(554), .Q_N(3000), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5140  (.CLK(clk_cts_n0), .D(2522), .Q(552), .Q_N(3001), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5141  (.CLK(clk_cts_n0), .D(2525), .Q(453), .Q_N(3002), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5142  (.CLK(clk_cts_n0), .D(2528), .Q(454), .Q_N(3003), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5143  (.CLK(clk_cts_n0), .D(2531), .Q(2021), .Q_N(3004), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5144  (.CLK(clk_cts_n0), .D(2534), .Q(2014), .Q_N(3005), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5145  (.CLK(clk_cts_n0), .D(2538), .Q(2138), .Q_N(3006), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5146  (.CLK(clk_cts_n2), .D(2543), .Q(511), .Q_N(3007), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5151  (.CLK(clk_cts_n0), .D(2552), .Q(1523), .Q_N(3008), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5152  (.CLK(clk_cts_n6), .D(2555), .Q(1555), .Q_N(3009), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5153  (.CLK(clk_cts_n0), .D(2566), .Q(544), .Q_N(3010), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5154  (.CLK(clk_cts_n4), .D(2568), .Q(539), .Q_N(3011), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5155  (.CLK(clk_cts_n0), .D(2574), .Q(546), .Q_N(3012), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5156  (.CLK(clk_cts_n4), .D(2578), .Q(1886), .Q_N(2197), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5157  (.CLK(clk_cts_n0), .D(2584), .Q(1543), .Q_N(3013), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5158  (.CLK(clk_cts_n2), .D(2587), .Q(1525), .Q_N(3014), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5159  (.CLK(clk_cts_n0), .D(2591), .Q(1196), .Q_N(562), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5160  (.CLK(clk_cts_n2), .D(2597), .Q(1193), .Q_N(3015), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5161  (.CLK(clk_cts_n0), .D(2606), .Q(2175), .Q_N(3016), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5166  (.CLK(clk_cts_n0), .D(2629), .Q(481), .Q_N(3017), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5167  (.CLK(clk_cts_n0), .D(2667), .Q(675), .Q_N(3018), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5168  (.CLK(clk_cts_n0), .D(2685), .Q(721), .Q_N(3019), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5169  (.CLK(clk_cts_n0), .D(141), .Q(138), .Q_N(3020), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5170  (.CLK(clk_cts_n0), .D(166), .Q(142), .Q_N(3021), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5171  (.CLK(clk_cts_n0), .D(188), .Q(167), .Q_N(3022), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5172  (.CLK(clk_cts_n0), .D(210), .Q(189), .Q_N(3023), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5173  (.CLK(clk_cts_n2), .D(231), .Q(211), .Q_N(3024), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5174  (.CLK(clk_cts_n0), .D(252), .Q(232), .Q_N(3025), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5175  (.CLK(clk_cts_n2), .D(278), .Q(253), .Q_N(3026), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5176  (.CLK(clk_cts_n0), .D(302), .Q(279), .Q_N(3027), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5177  (.CLK(clk_cts_n6), .D(326), .Q(303), .Q_N(3028), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5178  (.CLK(clk_cts_n0), .D(348), .Q(327), .Q_N(3029), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5179  (.CLK(clk_cts_n6), .D(372), .Q(349), .Q_N(3030), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5180  (.CLK(clk_cts_n0), .D(395), .Q(373), .Q_N(3031), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5181  (.CLK(clk_cts_n4), .D(416), .Q(396), .Q_N(3032), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5182  (.CLK(clk_cts_n0), .D(437), .Q(417), .Q_N(3033), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5183  (.CLK(clk_cts_n2), .D(1998), .Q(1995), .Q_N(2672), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5189  (.CLK(clk_cts_n0), .D(256), .Q(2214), .Q_N(3034), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5190  (.CLK(clk_cts_n2), .D(281), .Q(2231), .Q_N(3035), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5191  (.CLK(clk_cts_n0), .D(305), .Q(2250), .Q_N(3036), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5192  (.CLK(clk_cts_n2), .D(329), .Q(2269), .Q_N(3037), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5193  (.CLK(clk_cts_n3), .D(352), .Q(2294), .Q_N(3038), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5194  (.CLK(clk_cts_n3), .D(375), .Q(2310), .Q_N(3039), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5195  (.CLK(clk_cts_n3), .D(398), .Q(2329), .Q_N(3040), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5196  (.CLK(clk_cts_n3), .D(419), .Q(2347), .Q_N(3041), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5197  (.CLK(clk_cts_n3), .D(442), .Q(438), .Q_N(1238), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5198  (.CLK(clk_cts_n3), .D(447), .Q(443), .Q_N(1232), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5199  (.CLK(clk_cts_n9), .D(452), .Q(448), .Q_N(2148), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5200  (.CLK(clk_cts_n3), .D(2008), .Q(2000), .Q_N(3042), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5201  (.CLK(clk_cts_n9), .D(480), .Q(474), .Q_N(3043), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5202  (.CLK(clk_cts_n3), .D(507), .Q(2121), .Q_N(1249), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5203  (.CLK(clk_cts_n9), .D(2030), .Q(2009), .Q_N(2467), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5204  (.CLK(clk_cts_n3), .D(538), .Q(531), .Q_N(1235), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5205  (.CLK(clk_cts_n9), .D(582), .Q(577), .Q_N(1230), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5206  (.CLK(clk_cts_n0), .D(586), .Q(583), .Q_N(3044), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5207  (.CLK(clk_cts_n6), .D(704), .Q(678), .Q_N(3045), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5208  (.CLK(clk_cts_n0), .D(735), .Q(724), .Q_N(3046), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5209  (.CLK(clk_cts_n6), .D(765), .Q(753), .Q_N(3047), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5210  (.CLK(clk_cts_n0), .D(794), .Q(152), .Q_N(3048), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5211  (.CLK(clk_cts_n4), .D(823), .Q(175), .Q_N(3049), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5212  (.CLK(clk_cts_n0), .D(852), .Q(194), .Q_N(3050), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5213  (.CLK(clk_cts_n4), .D(881), .Q(218), .Q_N(3051), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5214  (.CLK(clk_cts_n0), .D(908), .Q(239), .Q_N(3052), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5215  (.CLK(clk_cts_n2), .D(2133), .Q(3053), .Q_N(2196), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5216  (.CLK(clk_cts_n0), .D(921), .Q(258), .Q_N(3054), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5217  (.CLK(clk_cts_n2), .D(932), .Q(283), .Q_N(3055), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5218  (.CLK(clk_cts_n3), .D(943), .Q(307), .Q_N(3056), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5219  (.CLK(clk_cts_n9), .D(954), .Q(331), .Q_N(3057), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5220  (.CLK(clk_cts_n3), .D(965), .Q(355), .Q_N(3058), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5221  (.CLK(clk_cts_n3), .D(976), .Q(378), .Q_N(3059), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5222  (.CLK(clk_cts_n3), .D(989), .Q(400), .Q_N(3060), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5223  (.CLK(clk_cts_n3), .D(1000), .Q(421), .Q_N(3061), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5224  (.CLK(clk_cts_n3), .D(1008), .Q(1006), .Q_N(3062), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5225  (.CLK(clk_cts_n3), .D(1012), .Q(1010), .Q_N(3063), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5226  (.CLK(clk_cts_n3), .D(1017), .Q(1013), .Q_N(3064), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5227  (.CLK(clk_cts_n3), .D(1021), .Q(1019), .Q_N(3065), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5228  (.CLK(clk_cts_n10), .D(1025), .Q(1023), .Q_N(3066), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5229  (.CLK(clk_cts_n3), .D(1030), .Q(1026), .Q_N(3067), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5230  (.CLK(clk_cts_n10), .D(1035), .Q(1031), .Q_N(3068), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5231  (.CLK(clk_cts_n3), .D(1039), .Q(1036), .Q_N(3069), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5232  (.CLK(clk_cts_n10), .D(1218), .Q(1216), .Q_N(2158), .RESET_B(3), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5233  (.CLK(clk_cts_n3), .D(1291), .Q(1288), .Q_N(2150), .RESET_B(3), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5234  (.CLK(clk_cts_n9), .D(1318), .Q(1316), .Q_N(2159), .RESET_B(3), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5235  (.CLK(clk_cts_n0), .D(1348), .Q(1346), .Q_N(2152), .RESET_B(2694), .SET_B(3));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5236  (.CLK(clk_cts_n6), .D(1370), .Q(1368), .Q_N(2155), .RESET_B(3), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$5237  (.CLK(clk_cts_n0), .D(1385), .Q(1383), .Q_N(2149), .RESET_B(3), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8804  (.CLK(clk_cts_n6), .D(1409), .Q(1386), .Q_N(3070), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8805  (.CLK(clk_cts_n0), .D(1421), .Q(1410), .Q_N(3071), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8806  (.CLK(clk_cts_n4), .D(1444), .Q(2147), .Q_N(3072), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8807  (.CLK(clk_cts_n0), .D(1452), .Q(1449), .Q_N(3073), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8808  (.CLK(clk_cts_n4), .D(1472), .Q(1453), .Q_N(3074), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8809  (.CLK(clk_cts_n0), .D(1490), .Q(1488), .Q_N(3075), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8810  (.CLK(clk_cts_n2), .D(1503), .Q(1491), .Q_N(3076), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\$auto$ff.cc:266:slice$8811  (.CLK(clk_cts_n0), .D(1512), .Q(1504), .Q_N(3077), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7456  (.CLK(clk_cts_n2), .D(1653), .Q(1513), .Q_N(3078), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7679  (.CLK(clk_cts_n3), .D(1922), .Q(234), .Q_N(3079), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7680  (.CLK(clk_cts_n9), .D(1926), .Q(1923), .Q_N(2199), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7681  (.CLK(clk_cts_n3), .D(1932), .Q(516), .Q_N(3080), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7682  (.CLK(clk_cts_n9), .D(1936), .Q(286), .Q_N(3081), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7683  (.CLK(clk_cts_n3), .D(1940), .Q(518), .Q_N(3082), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7684  (.CLK(clk_cts_n3), .D(1944), .Q(145), .Q_N(3083), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7685  (.CLK(clk_cts_n3), .D(1950), .Q(169), .Q_N(3084), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7686  (.CLK(clk_cts_n3), .D(1956), .Q(191), .Q_N(3085), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7687  (.CLK(clk_cts_n3), .D(1962), .Q(213), .Q_N(3086), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7689  (.CLK(clk_cts_n3), .D(1966), .Q(1963), .Q_N(3087), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__dfbbp_1 \$flatten \CPU.\ALU.\$auto$ff.cc:266:slice$7690  (.CLK(clk_cts_n3), .D(1982), .Q(550), .Q_N(2279), .RESET_B(2694), .SET_B(2694));
  sky130_fd_sc_hd__conb_1 conb_T0Y0 (.HI(tie_high_T0Y0), .LO(tie_low_T0Y0));
  sky130_fd_sc_hd__conb_1 conb_T0Y1 (.HI(tie_high_T0Y1), .LO(tie_low_T0Y1));
  sky130_fd_sc_hd__conb_1 conb_T0Y10 (.HI(tie_high_T0Y10), .LO(tie_low_T0Y10));
  sky130_fd_sc_hd__conb_1 conb_T0Y11 (.HI(tie_high_T0Y11), .LO(tie_low_T0Y11));
  sky130_fd_sc_hd__conb_1 conb_T0Y12 (.HI(tie_high_T0Y12), .LO(tie_low_T0Y12));
  sky130_fd_sc_hd__conb_1 conb_T0Y13 (.HI(tie_high_T0Y13), .LO(tie_low_T0Y13));
  sky130_fd_sc_hd__conb_1 conb_T0Y14 (.HI(tie_high_T0Y14), .LO(tie_low_T0Y14));
  sky130_fd_sc_hd__conb_1 conb_T0Y15 (.HI(tie_high_T0Y15), .LO(tie_low_T0Y15));
  sky130_fd_sc_hd__conb_1 conb_T0Y16 (.HI(tie_high_T0Y16), .LO(tie_low_T0Y16));
  sky130_fd_sc_hd__conb_1 conb_T0Y17 (.HI(tie_high_T0Y17), .LO(tie_low_T0Y17));
  sky130_fd_sc_hd__conb_1 conb_T0Y18 (.HI(tie_high_T0Y18), .LO(tie_low_T0Y18));
  sky130_fd_sc_hd__conb_1 conb_T0Y19 (.HI(tie_high_T0Y19), .LO(tie_low_T0Y19));
  sky130_fd_sc_hd__conb_1 conb_T0Y2 (.HI(tie_high_T0Y2), .LO(tie_low_T0Y2));
  sky130_fd_sc_hd__conb_1 conb_T0Y20 (.HI(tie_high_T0Y20), .LO(tie_low_T0Y20));
  sky130_fd_sc_hd__conb_1 conb_T0Y21 (.HI(tie_high_T0Y21), .LO(tie_low_T0Y21));
  sky130_fd_sc_hd__conb_1 conb_T0Y22 (.HI(tie_high_T0Y22), .LO(tie_low_T0Y22));
  sky130_fd_sc_hd__conb_1 conb_T0Y23 (.HI(tie_high_T0Y23), .LO(tie_low_T0Y23));
  sky130_fd_sc_hd__conb_1 conb_T0Y24 (.HI(tie_high_T0Y24), .LO(tie_low_T0Y24));
  sky130_fd_sc_hd__conb_1 conb_T0Y25 (.HI(tie_high_T0Y25), .LO(tie_low_T0Y25));
  sky130_fd_sc_hd__conb_1 conb_T0Y26 (.HI(tie_high_T0Y26), .LO(tie_low_T0Y26));
  sky130_fd_sc_hd__conb_1 conb_T0Y27 (.HI(tie_high_T0Y27), .LO(tie_low_T0Y27));
  sky130_fd_sc_hd__conb_1 conb_T0Y28 (.HI(tie_high_T0Y28), .LO(tie_low_T0Y28));
  sky130_fd_sc_hd__conb_1 conb_T0Y29 (.HI(tie_high_T0Y29), .LO(tie_low_T0Y29));
  sky130_fd_sc_hd__conb_1 conb_T0Y3 (.HI(tie_high_T0Y3), .LO(tie_low_T0Y3));
  sky130_fd_sc_hd__conb_1 conb_T0Y30 (.HI(tie_high_T0Y30), .LO(tie_low_T0Y30));
  sky130_fd_sc_hd__conb_1 conb_T0Y31 (.HI(tie_high_T0Y31), .LO(tie_low_T0Y31));
  sky130_fd_sc_hd__conb_1 conb_T0Y32 (.HI(tie_high_T0Y32), .LO(tie_low_T0Y32));
  sky130_fd_sc_hd__conb_1 conb_T0Y33 (.HI(tie_high_T0Y33), .LO(tie_low_T0Y33));
  sky130_fd_sc_hd__conb_1 conb_T0Y34 (.HI(tie_high_T0Y34), .LO(tie_low_T0Y34));
  sky130_fd_sc_hd__conb_1 conb_T0Y35 (.HI(tie_high_T0Y35), .LO(tie_low_T0Y35));
  sky130_fd_sc_hd__conb_1 conb_T0Y36 (.HI(tie_high_T0Y36), .LO(tie_low_T0Y36));
  sky130_fd_sc_hd__conb_1 conb_T0Y37 (.HI(tie_high_T0Y37), .LO(tie_low_T0Y37));
  sky130_fd_sc_hd__conb_1 conb_T0Y38 (.HI(tie_high_T0Y38), .LO(tie_low_T0Y38));
  sky130_fd_sc_hd__conb_1 conb_T0Y39 (.HI(tie_high_T0Y39), .LO(tie_low_T0Y39));
  sky130_fd_sc_hd__conb_1 conb_T0Y4 (.HI(tie_high_T0Y4), .LO(tie_low_T0Y4));
  sky130_fd_sc_hd__conb_1 conb_T0Y40 (.HI(tie_high_T0Y40), .LO(tie_low_T0Y40));
  sky130_fd_sc_hd__conb_1 conb_T0Y41 (.HI(tie_high_T0Y41), .LO(tie_low_T0Y41));
  sky130_fd_sc_hd__conb_1 conb_T0Y42 (.HI(tie_high_T0Y42), .LO(tie_low_T0Y42));
  sky130_fd_sc_hd__conb_1 conb_T0Y43 (.HI(tie_high_T0Y43), .LO(tie_low_T0Y43));
  sky130_fd_sc_hd__conb_1 conb_T0Y44 (.HI(tie_high_T0Y44), .LO(tie_low_T0Y44));
  sky130_fd_sc_hd__conb_1 conb_T0Y45 (.HI(tie_high_T0Y45), .LO(tie_low_T0Y45));
  sky130_fd_sc_hd__conb_1 conb_T0Y46 (.HI(tie_high_T0Y46), .LO(tie_low_T0Y46));
  sky130_fd_sc_hd__conb_1 conb_T0Y47 (.HI(tie_high_T0Y47), .LO(tie_low_T0Y47));
  sky130_fd_sc_hd__conb_1 conb_T0Y48 (.HI(tie_high_T0Y48), .LO(tie_low_T0Y48));
  sky130_fd_sc_hd__conb_1 conb_T0Y49 (.HI(tie_high_T0Y49), .LO(tie_low_T0Y49));
  sky130_fd_sc_hd__conb_1 conb_T0Y5 (.HI(tie_high_T0Y5), .LO(tie_low_T0Y5));
  sky130_fd_sc_hd__conb_1 conb_T0Y50 (.HI(tie_high_T0Y50), .LO(tie_low_T0Y50));
  sky130_fd_sc_hd__conb_1 conb_T0Y51 (.HI(tie_high_T0Y51), .LO(tie_low_T0Y51));
  sky130_fd_sc_hd__conb_1 conb_T0Y52 (.HI(tie_high_T0Y52), .LO(tie_low_T0Y52));
  sky130_fd_sc_hd__conb_1 conb_T0Y53 (.HI(tie_high_T0Y53), .LO(tie_low_T0Y53));
  sky130_fd_sc_hd__conb_1 conb_T0Y54 (.HI(tie_high_T0Y54), .LO(tie_low_T0Y54));
  sky130_fd_sc_hd__conb_1 conb_T0Y55 (.HI(tie_high_T0Y55), .LO(tie_low_T0Y55));
  sky130_fd_sc_hd__conb_1 conb_T0Y56 (.HI(tie_high_T0Y56), .LO(tie_low_T0Y56));
  sky130_fd_sc_hd__conb_1 conb_T0Y57 (.HI(tie_high_T0Y57), .LO(tie_low_T0Y57));
  sky130_fd_sc_hd__conb_1 conb_T0Y58 (.HI(tie_high_T0Y58), .LO(tie_low_T0Y58));
  sky130_fd_sc_hd__conb_1 conb_T0Y59 (.HI(tie_high_T0Y59), .LO(tie_low_T0Y59));
  sky130_fd_sc_hd__conb_1 conb_T0Y6 (.HI(tie_high_T0Y6), .LO(tie_low_T0Y6));
  sky130_fd_sc_hd__conb_1 conb_T0Y60 (.HI(tie_high_T0Y60), .LO(tie_low_T0Y60));
  sky130_fd_sc_hd__conb_1 conb_T0Y61 (.HI(tie_high_T0Y61), .LO(tie_low_T0Y61));
  sky130_fd_sc_hd__conb_1 conb_T0Y62 (.HI(tie_high_T0Y62), .LO(tie_low_T0Y62));
  sky130_fd_sc_hd__conb_1 conb_T0Y63 (.HI(tie_high_T0Y63), .LO(tie_low_T0Y63));
  sky130_fd_sc_hd__conb_1 conb_T0Y64 (.HI(tie_high_T0Y64), .LO(tie_low_T0Y64));
  sky130_fd_sc_hd__conb_1 conb_T0Y65 (.HI(tie_high_T0Y65), .LO(tie_low_T0Y65));
  sky130_fd_sc_hd__conb_1 conb_T0Y66 (.HI(tie_high_T0Y66), .LO(tie_low_T0Y66));
  sky130_fd_sc_hd__conb_1 conb_T0Y67 (.HI(tie_high_T0Y67), .LO(tie_low_T0Y67));
  sky130_fd_sc_hd__conb_1 conb_T0Y68 (.HI(tie_high_T0Y68), .LO(tie_low_T0Y68));
  sky130_fd_sc_hd__conb_1 conb_T0Y69 (.HI(tie_high_T0Y69), .LO(tie_low_T0Y69));
  sky130_fd_sc_hd__conb_1 conb_T0Y7 (.HI(tie_high_T0Y7), .LO(tie_low_T0Y7));
  sky130_fd_sc_hd__conb_1 conb_T0Y70 (.HI(tie_high_T0Y70), .LO(tie_low_T0Y70));
  sky130_fd_sc_hd__conb_1 conb_T0Y71 (.HI(tie_high_T0Y71), .LO(tie_low_T0Y71));
  sky130_fd_sc_hd__conb_1 conb_T0Y72 (.HI(tie_high_T0Y72), .LO(tie_low_T0Y72));
  sky130_fd_sc_hd__conb_1 conb_T0Y73 (.HI(tie_high_T0Y73), .LO(tie_low_T0Y73));
  sky130_fd_sc_hd__conb_1 conb_T0Y74 (.HI(tie_high_T0Y74), .LO(tie_low_T0Y74));
  sky130_fd_sc_hd__conb_1 conb_T0Y75 (.HI(tie_high_T0Y75), .LO(tie_low_T0Y75));
  sky130_fd_sc_hd__conb_1 conb_T0Y76 (.HI(tie_high_T0Y76), .LO(tie_low_T0Y76));
  sky130_fd_sc_hd__conb_1 conb_T0Y77 (.HI(tie_high_T0Y77), .LO(tie_low_T0Y77));
  sky130_fd_sc_hd__conb_1 conb_T0Y78 (.HI(tie_high_T0Y78), .LO(tie_low_T0Y78));
  sky130_fd_sc_hd__conb_1 conb_T0Y79 (.HI(tie_high_T0Y79), .LO(tie_low_T0Y79));
  sky130_fd_sc_hd__conb_1 conb_T0Y8 (.HI(tie_high_T0Y8), .LO(tie_low_T0Y8));
  sky130_fd_sc_hd__conb_1 conb_T0Y80 (.HI(tie_high_T0Y80), .LO(tie_low_T0Y80));
  sky130_fd_sc_hd__conb_1 conb_T0Y81 (.HI(tie_high_T0Y81), .LO(tie_low_T0Y81));
  sky130_fd_sc_hd__conb_1 conb_T0Y82 (.HI(tie_high_T0Y82), .LO(tie_low_T0Y82));
  sky130_fd_sc_hd__conb_1 conb_T0Y83 (.HI(tie_high_T0Y83), .LO(tie_low_T0Y83));
  sky130_fd_sc_hd__conb_1 conb_T0Y84 (.HI(tie_high_T0Y84), .LO(tie_low_T0Y84));
  sky130_fd_sc_hd__conb_1 conb_T0Y85 (.HI(tie_high_T0Y85), .LO(tie_low_T0Y85));
  sky130_fd_sc_hd__conb_1 conb_T0Y86 (.HI(tie_high_T0Y86), .LO(tie_low_T0Y86));
  sky130_fd_sc_hd__conb_1 conb_T0Y87 (.HI(tie_high_T0Y87), .LO(tie_low_T0Y87));
  sky130_fd_sc_hd__conb_1 conb_T0Y88 (.HI(tie_high_T0Y88), .LO(tie_low_T0Y88));
  sky130_fd_sc_hd__conb_1 conb_T0Y89 (.HI(tie_high_T0Y89), .LO(tie_low_T0Y89));
  sky130_fd_sc_hd__conb_1 conb_T0Y9 (.HI(tie_high_T0Y9), .LO(tie_low_T0Y9));
  sky130_fd_sc_hd__conb_1 conb_T10Y0 (.HI(tie_high_T10Y0), .LO(tie_low_T10Y0));
  sky130_fd_sc_hd__conb_1 conb_T10Y1 (.HI(tie_high_T10Y1), .LO(tie_low_T10Y1));
  sky130_fd_sc_hd__conb_1 conb_T10Y10 (.HI(tie_high_T10Y10), .LO(tie_low_T10Y10));
  sky130_fd_sc_hd__conb_1 conb_T10Y11 (.HI(tie_high_T10Y11), .LO(tie_low_T10Y11));
  sky130_fd_sc_hd__conb_1 conb_T10Y12 (.HI(tie_high_T10Y12), .LO(tie_low_T10Y12));
  sky130_fd_sc_hd__conb_1 conb_T10Y13 (.HI(tie_high_T10Y13), .LO(tie_low_T10Y13));
  sky130_fd_sc_hd__conb_1 conb_T10Y14 (.HI(tie_high_T10Y14), .LO(tie_low_T10Y14));
  sky130_fd_sc_hd__conb_1 conb_T10Y15 (.HI(tie_high_T10Y15), .LO(tie_low_T10Y15));
  sky130_fd_sc_hd__conb_1 conb_T10Y16 (.HI(tie_high_T10Y16), .LO(tie_low_T10Y16));
  sky130_fd_sc_hd__conb_1 conb_T10Y17 (.HI(tie_high_T10Y17), .LO(tie_low_T10Y17));
  sky130_fd_sc_hd__conb_1 conb_T10Y18 (.HI(tie_high_T10Y18), .LO(tie_low_T10Y18));
  sky130_fd_sc_hd__conb_1 conb_T10Y19 (.HI(tie_high_T10Y19), .LO(tie_low_T10Y19));
  sky130_fd_sc_hd__conb_1 conb_T10Y2 (.HI(tie_high_T10Y2), .LO(tie_low_T10Y2));
  sky130_fd_sc_hd__conb_1 conb_T10Y20 (.HI(tie_high_T10Y20), .LO(tie_low_T10Y20));
  sky130_fd_sc_hd__conb_1 conb_T10Y21 (.HI(tie_high_T10Y21), .LO(tie_low_T10Y21));
  sky130_fd_sc_hd__conb_1 conb_T10Y22 (.HI(tie_high_T10Y22), .LO(tie_low_T10Y22));
  sky130_fd_sc_hd__conb_1 conb_T10Y23 (.HI(tie_high_T10Y23), .LO(tie_low_T10Y23));
  sky130_fd_sc_hd__conb_1 conb_T10Y24 (.HI(tie_high_T10Y24), .LO(tie_low_T10Y24));
  sky130_fd_sc_hd__conb_1 conb_T10Y25 (.HI(tie_high_T10Y25), .LO(tie_low_T10Y25));
  sky130_fd_sc_hd__conb_1 conb_T10Y26 (.HI(tie_high_T10Y26), .LO(tie_low_T10Y26));
  sky130_fd_sc_hd__conb_1 conb_T10Y27 (.HI(tie_high_T10Y27), .LO(tie_low_T10Y27));
  sky130_fd_sc_hd__conb_1 conb_T10Y28 (.HI(tie_high_T10Y28), .LO(tie_low_T10Y28));
  sky130_fd_sc_hd__conb_1 conb_T10Y29 (.HI(tie_high_T10Y29), .LO(tie_low_T10Y29));
  sky130_fd_sc_hd__conb_1 conb_T10Y3 (.HI(tie_high_T10Y3), .LO(tie_low_T10Y3));
  sky130_fd_sc_hd__conb_1 conb_T10Y30 (.HI(tie_high_T10Y30), .LO(tie_low_T10Y30));
  sky130_fd_sc_hd__conb_1 conb_T10Y31 (.HI(tie_high_T10Y31), .LO(tie_low_T10Y31));
  sky130_fd_sc_hd__conb_1 conb_T10Y32 (.HI(tie_high_T10Y32), .LO(tie_low_T10Y32));
  sky130_fd_sc_hd__conb_1 conb_T10Y33 (.HI(tie_high_T10Y33), .LO(tie_low_T10Y33));
  sky130_fd_sc_hd__conb_1 conb_T10Y34 (.HI(tie_high_T10Y34), .LO(tie_low_T10Y34));
  sky130_fd_sc_hd__conb_1 conb_T10Y35 (.HI(tie_high_T10Y35), .LO(tie_low_T10Y35));
  sky130_fd_sc_hd__conb_1 conb_T10Y36 (.HI(tie_high_T10Y36), .LO(tie_low_T10Y36));
  sky130_fd_sc_hd__conb_1 conb_T10Y37 (.HI(tie_high_T10Y37), .LO(tie_low_T10Y37));
  sky130_fd_sc_hd__conb_1 conb_T10Y38 (.HI(tie_high_T10Y38), .LO(tie_low_T10Y38));
  sky130_fd_sc_hd__conb_1 conb_T10Y39 (.HI(tie_high_T10Y39), .LO(tie_low_T10Y39));
  sky130_fd_sc_hd__conb_1 conb_T10Y4 (.HI(tie_high_T10Y4), .LO(tie_low_T10Y4));
  sky130_fd_sc_hd__conb_1 conb_T10Y40 (.HI(tie_high_T10Y40), .LO(tie_low_T10Y40));
  sky130_fd_sc_hd__conb_1 conb_T10Y41 (.HI(tie_high_T10Y41), .LO(tie_low_T10Y41));
  sky130_fd_sc_hd__conb_1 conb_T10Y42 (.HI(tie_high_T10Y42), .LO(tie_low_T10Y42));
  sky130_fd_sc_hd__conb_1 conb_T10Y43 (.HI(tie_high_T10Y43), .LO(tie_low_T10Y43));
  sky130_fd_sc_hd__conb_1 conb_T10Y44 (.HI(tie_high_T10Y44), .LO(tie_low_T10Y44));
  sky130_fd_sc_hd__conb_1 conb_T10Y45 (.HI(tie_high_T10Y45), .LO(tie_low_T10Y45));
  sky130_fd_sc_hd__conb_1 conb_T10Y46 (.HI(tie_high_T10Y46), .LO(tie_low_T10Y46));
  sky130_fd_sc_hd__conb_1 conb_T10Y47 (.HI(tie_high_T10Y47), .LO(tie_low_T10Y47));
  sky130_fd_sc_hd__conb_1 conb_T10Y48 (.HI(tie_high_T10Y48), .LO(tie_low_T10Y48));
  sky130_fd_sc_hd__conb_1 conb_T10Y49 (.HI(tie_high_T10Y49), .LO(tie_low_T10Y49));
  sky130_fd_sc_hd__conb_1 conb_T10Y5 (.HI(tie_high_T10Y5), .LO(tie_low_T10Y5));
  sky130_fd_sc_hd__conb_1 conb_T10Y50 (.HI(tie_high_T10Y50), .LO(tie_low_T10Y50));
  sky130_fd_sc_hd__conb_1 conb_T10Y51 (.HI(tie_high_T10Y51), .LO(tie_low_T10Y51));
  sky130_fd_sc_hd__conb_1 conb_T10Y52 (.HI(tie_high_T10Y52), .LO(tie_low_T10Y52));
  sky130_fd_sc_hd__conb_1 conb_T10Y53 (.HI(tie_high_T10Y53), .LO(tie_low_T10Y53));
  sky130_fd_sc_hd__conb_1 conb_T10Y54 (.HI(tie_high_T10Y54), .LO(tie_low_T10Y54));
  sky130_fd_sc_hd__conb_1 conb_T10Y55 (.HI(tie_high_T10Y55), .LO(tie_low_T10Y55));
  sky130_fd_sc_hd__conb_1 conb_T10Y56 (.HI(tie_high_T10Y56), .LO(tie_low_T10Y56));
  sky130_fd_sc_hd__conb_1 conb_T10Y57 (.HI(tie_high_T10Y57), .LO(tie_low_T10Y57));
  sky130_fd_sc_hd__conb_1 conb_T10Y58 (.HI(tie_high_T10Y58), .LO(tie_low_T10Y58));
  sky130_fd_sc_hd__conb_1 conb_T10Y59 (.HI(tie_high_T10Y59), .LO(tie_low_T10Y59));
  sky130_fd_sc_hd__conb_1 conb_T10Y6 (.HI(tie_high_T10Y6), .LO(tie_low_T10Y6));
  sky130_fd_sc_hd__conb_1 conb_T10Y60 (.HI(tie_high_T10Y60), .LO(tie_low_T10Y60));
  sky130_fd_sc_hd__conb_1 conb_T10Y61 (.HI(tie_high_T10Y61), .LO(tie_low_T10Y61));
  sky130_fd_sc_hd__conb_1 conb_T10Y62 (.HI(tie_high_T10Y62), .LO(tie_low_T10Y62));
  sky130_fd_sc_hd__conb_1 conb_T10Y63 (.HI(tie_high_T10Y63), .LO(tie_low_T10Y63));
  sky130_fd_sc_hd__conb_1 conb_T10Y64 (.HI(tie_high_T10Y64), .LO(tie_low_T10Y64));
  sky130_fd_sc_hd__conb_1 conb_T10Y65 (.HI(tie_high_T10Y65), .LO(tie_low_T10Y65));
  sky130_fd_sc_hd__conb_1 conb_T10Y66 (.HI(tie_high_T10Y66), .LO(tie_low_T10Y66));
  sky130_fd_sc_hd__conb_1 conb_T10Y67 (.HI(tie_high_T10Y67), .LO(tie_low_T10Y67));
  sky130_fd_sc_hd__conb_1 conb_T10Y68 (.HI(tie_high_T10Y68), .LO(tie_low_T10Y68));
  sky130_fd_sc_hd__conb_1 conb_T10Y69 (.HI(tie_high_T10Y69), .LO(tie_low_T10Y69));
  sky130_fd_sc_hd__conb_1 conb_T10Y7 (.HI(tie_high_T10Y7), .LO(tie_low_T10Y7));
  sky130_fd_sc_hd__conb_1 conb_T10Y70 (.HI(tie_high_T10Y70), .LO(tie_low_T10Y70));
  sky130_fd_sc_hd__conb_1 conb_T10Y71 (.HI(tie_high_T10Y71), .LO(tie_low_T10Y71));
  sky130_fd_sc_hd__conb_1 conb_T10Y72 (.HI(tie_high_T10Y72), .LO(tie_low_T10Y72));
  sky130_fd_sc_hd__conb_1 conb_T10Y73 (.HI(tie_high_T10Y73), .LO(tie_low_T10Y73));
  sky130_fd_sc_hd__conb_1 conb_T10Y74 (.HI(tie_high_T10Y74), .LO(tie_low_T10Y74));
  sky130_fd_sc_hd__conb_1 conb_T10Y75 (.HI(tie_high_T10Y75), .LO(tie_low_T10Y75));
  sky130_fd_sc_hd__conb_1 conb_T10Y76 (.HI(tie_high_T10Y76), .LO(tie_low_T10Y76));
  sky130_fd_sc_hd__conb_1 conb_T10Y77 (.HI(tie_high_T10Y77), .LO(tie_low_T10Y77));
  sky130_fd_sc_hd__conb_1 conb_T10Y78 (.HI(tie_high_T10Y78), .LO(tie_low_T10Y78));
  sky130_fd_sc_hd__conb_1 conb_T10Y79 (.HI(tie_high_T10Y79), .LO(tie_low_T10Y79));
  sky130_fd_sc_hd__conb_1 conb_T10Y8 (.HI(tie_high_T10Y8), .LO(tie_low_T10Y8));
  sky130_fd_sc_hd__conb_1 conb_T10Y80 (.HI(tie_high_T10Y80), .LO(tie_low_T10Y80));
  sky130_fd_sc_hd__conb_1 conb_T10Y81 (.HI(tie_high_T10Y81), .LO(tie_low_T10Y81));
  sky130_fd_sc_hd__conb_1 conb_T10Y82 (.HI(tie_high_T10Y82), .LO(tie_low_T10Y82));
  sky130_fd_sc_hd__conb_1 conb_T10Y83 (.HI(tie_high_T10Y83), .LO(tie_low_T10Y83));
  sky130_fd_sc_hd__conb_1 conb_T10Y84 (.HI(tie_high_T10Y84), .LO(tie_low_T10Y84));
  sky130_fd_sc_hd__conb_1 conb_T10Y85 (.HI(tie_high_T10Y85), .LO(tie_low_T10Y85));
  sky130_fd_sc_hd__conb_1 conb_T10Y86 (.HI(tie_high_T10Y86), .LO(tie_low_T10Y86));
  sky130_fd_sc_hd__conb_1 conb_T10Y87 (.HI(tie_high_T10Y87), .LO(tie_low_T10Y87));
  sky130_fd_sc_hd__conb_1 conb_T10Y88 (.HI(tie_high_T10Y88), .LO(tie_low_T10Y88));
  sky130_fd_sc_hd__conb_1 conb_T10Y89 (.HI(tie_high_T10Y89), .LO(tie_low_T10Y89));
  sky130_fd_sc_hd__conb_1 conb_T10Y9 (.HI(tie_high_T10Y9), .LO(tie_low_T10Y9));
  sky130_fd_sc_hd__conb_1 conb_T11Y0 (.HI(tie_high_T11Y0), .LO(tie_low_T11Y0));
  sky130_fd_sc_hd__conb_1 conb_T11Y1 (.HI(tie_high_T11Y1), .LO(tie_low_T11Y1));
  sky130_fd_sc_hd__conb_1 conb_T11Y10 (.HI(tie_high_T11Y10), .LO(tie_low_T11Y10));
  sky130_fd_sc_hd__conb_1 conb_T11Y11 (.HI(tie_high_T11Y11), .LO(tie_low_T11Y11));
  sky130_fd_sc_hd__conb_1 conb_T11Y12 (.HI(tie_high_T11Y12), .LO(tie_low_T11Y12));
  sky130_fd_sc_hd__conb_1 conb_T11Y13 (.HI(tie_high_T11Y13), .LO(tie_low_T11Y13));
  sky130_fd_sc_hd__conb_1 conb_T11Y14 (.HI(tie_high_T11Y14), .LO(tie_low_T11Y14));
  sky130_fd_sc_hd__conb_1 conb_T11Y15 (.HI(tie_high_T11Y15), .LO(tie_low_T11Y15));
  sky130_fd_sc_hd__conb_1 conb_T11Y16 (.HI(tie_high_T11Y16), .LO(tie_low_T11Y16));
  sky130_fd_sc_hd__conb_1 conb_T11Y17 (.HI(tie_high_T11Y17), .LO(tie_low_T11Y17));
  sky130_fd_sc_hd__conb_1 conb_T11Y18 (.HI(tie_high_T11Y18), .LO(tie_low_T11Y18));
  sky130_fd_sc_hd__conb_1 conb_T11Y19 (.HI(tie_high_T11Y19), .LO(tie_low_T11Y19));
  sky130_fd_sc_hd__conb_1 conb_T11Y2 (.HI(tie_high_T11Y2), .LO(tie_low_T11Y2));
  sky130_fd_sc_hd__conb_1 conb_T11Y20 (.HI(tie_high_T11Y20), .LO(tie_low_T11Y20));
  sky130_fd_sc_hd__conb_1 conb_T11Y21 (.HI(tie_high_T11Y21), .LO(tie_low_T11Y21));
  sky130_fd_sc_hd__conb_1 conb_T11Y22 (.HI(tie_high_T11Y22), .LO(tie_low_T11Y22));
  sky130_fd_sc_hd__conb_1 conb_T11Y23 (.HI(tie_high_T11Y23), .LO(tie_low_T11Y23));
  sky130_fd_sc_hd__conb_1 conb_T11Y24 (.HI(tie_high_T11Y24), .LO(tie_low_T11Y24));
  sky130_fd_sc_hd__conb_1 conb_T11Y25 (.HI(tie_high_T11Y25), .LO(tie_low_T11Y25));
  sky130_fd_sc_hd__conb_1 conb_T11Y26 (.HI(tie_high_T11Y26), .LO(tie_low_T11Y26));
  sky130_fd_sc_hd__conb_1 conb_T11Y27 (.HI(tie_high_T11Y27), .LO(tie_low_T11Y27));
  sky130_fd_sc_hd__conb_1 conb_T11Y28 (.HI(tie_high_T11Y28), .LO(tie_low_T11Y28));
  sky130_fd_sc_hd__conb_1 conb_T11Y29 (.HI(tie_high_T11Y29), .LO(tie_low_T11Y29));
  sky130_fd_sc_hd__conb_1 conb_T11Y3 (.HI(tie_high_T11Y3), .LO(tie_low_T11Y3));
  sky130_fd_sc_hd__conb_1 conb_T11Y30 (.HI(tie_high_T11Y30), .LO(tie_low_T11Y30));
  sky130_fd_sc_hd__conb_1 conb_T11Y31 (.HI(tie_high_T11Y31), .LO(tie_low_T11Y31));
  sky130_fd_sc_hd__conb_1 conb_T11Y32 (.HI(tie_high_T11Y32), .LO(tie_low_T11Y32));
  sky130_fd_sc_hd__conb_1 conb_T11Y33 (.HI(tie_high_T11Y33), .LO(tie_low_T11Y33));
  sky130_fd_sc_hd__conb_1 conb_T11Y34 (.HI(tie_high_T11Y34), .LO(tie_low_T11Y34));
  sky130_fd_sc_hd__conb_1 conb_T11Y35 (.HI(tie_high_T11Y35), .LO(tie_low_T11Y35));
  sky130_fd_sc_hd__conb_1 conb_T11Y36 (.HI(tie_high_T11Y36), .LO(tie_low_T11Y36));
  sky130_fd_sc_hd__conb_1 conb_T11Y37 (.HI(tie_high_T11Y37), .LO(tie_low_T11Y37));
  sky130_fd_sc_hd__conb_1 conb_T11Y38 (.HI(tie_high_T11Y38), .LO(tie_low_T11Y38));
  sky130_fd_sc_hd__conb_1 conb_T11Y39 (.HI(tie_high_T11Y39), .LO(tie_low_T11Y39));
  sky130_fd_sc_hd__conb_1 conb_T11Y4 (.HI(tie_high_T11Y4), .LO(tie_low_T11Y4));
  sky130_fd_sc_hd__conb_1 conb_T11Y40 (.HI(tie_high_T11Y40), .LO(tie_low_T11Y40));
  sky130_fd_sc_hd__conb_1 conb_T11Y41 (.HI(tie_high_T11Y41), .LO(tie_low_T11Y41));
  sky130_fd_sc_hd__conb_1 conb_T11Y42 (.HI(tie_high_T11Y42), .LO(tie_low_T11Y42));
  sky130_fd_sc_hd__conb_1 conb_T11Y43 (.HI(tie_high_T11Y43), .LO(tie_low_T11Y43));
  sky130_fd_sc_hd__conb_1 conb_T11Y44 (.HI(tie_high_T11Y44), .LO(tie_low_T11Y44));
  sky130_fd_sc_hd__conb_1 conb_T11Y45 (.HI(tie_high_T11Y45), .LO(tie_low_T11Y45));
  sky130_fd_sc_hd__conb_1 conb_T11Y46 (.HI(tie_high_T11Y46), .LO(tie_low_T11Y46));
  sky130_fd_sc_hd__conb_1 conb_T11Y47 (.HI(tie_high_T11Y47), .LO(tie_low_T11Y47));
  sky130_fd_sc_hd__conb_1 conb_T11Y48 (.HI(tie_high_T11Y48), .LO(tie_low_T11Y48));
  sky130_fd_sc_hd__conb_1 conb_T11Y49 (.HI(tie_high_T11Y49), .LO(tie_low_T11Y49));
  sky130_fd_sc_hd__conb_1 conb_T11Y5 (.HI(tie_high_T11Y5), .LO(tie_low_T11Y5));
  sky130_fd_sc_hd__conb_1 conb_T11Y50 (.HI(tie_high_T11Y50), .LO(tie_low_T11Y50));
  sky130_fd_sc_hd__conb_1 conb_T11Y51 (.HI(tie_high_T11Y51), .LO(tie_low_T11Y51));
  sky130_fd_sc_hd__conb_1 conb_T11Y52 (.HI(tie_high_T11Y52), .LO(tie_low_T11Y52));
  sky130_fd_sc_hd__conb_1 conb_T11Y53 (.HI(tie_high_T11Y53), .LO(tie_low_T11Y53));
  sky130_fd_sc_hd__conb_1 conb_T11Y54 (.HI(tie_high_T11Y54), .LO(tie_low_T11Y54));
  sky130_fd_sc_hd__conb_1 conb_T11Y55 (.HI(tie_high_T11Y55), .LO(tie_low_T11Y55));
  sky130_fd_sc_hd__conb_1 conb_T11Y56 (.HI(tie_high_T11Y56), .LO(tie_low_T11Y56));
  sky130_fd_sc_hd__conb_1 conb_T11Y57 (.HI(tie_high_T11Y57), .LO(tie_low_T11Y57));
  sky130_fd_sc_hd__conb_1 conb_T11Y58 (.HI(tie_high_T11Y58), .LO(tie_low_T11Y58));
  sky130_fd_sc_hd__conb_1 conb_T11Y59 (.HI(tie_high_T11Y59), .LO(tie_low_T11Y59));
  sky130_fd_sc_hd__conb_1 conb_T11Y6 (.HI(tie_high_T11Y6), .LO(tie_low_T11Y6));
  sky130_fd_sc_hd__conb_1 conb_T11Y60 (.HI(tie_high_T11Y60), .LO(tie_low_T11Y60));
  sky130_fd_sc_hd__conb_1 conb_T11Y61 (.HI(tie_high_T11Y61), .LO(tie_low_T11Y61));
  sky130_fd_sc_hd__conb_1 conb_T11Y62 (.HI(tie_high_T11Y62), .LO(tie_low_T11Y62));
  sky130_fd_sc_hd__conb_1 conb_T11Y63 (.HI(tie_high_T11Y63), .LO(tie_low_T11Y63));
  sky130_fd_sc_hd__conb_1 conb_T11Y64 (.HI(tie_high_T11Y64), .LO(tie_low_T11Y64));
  sky130_fd_sc_hd__conb_1 conb_T11Y65 (.HI(tie_high_T11Y65), .LO(tie_low_T11Y65));
  sky130_fd_sc_hd__conb_1 conb_T11Y66 (.HI(tie_high_T11Y66), .LO(tie_low_T11Y66));
  sky130_fd_sc_hd__conb_1 conb_T11Y67 (.HI(tie_high_T11Y67), .LO(tie_low_T11Y67));
  sky130_fd_sc_hd__conb_1 conb_T11Y68 (.HI(tie_high_T11Y68), .LO(tie_low_T11Y68));
  sky130_fd_sc_hd__conb_1 conb_T11Y69 (.HI(tie_high_T11Y69), .LO(tie_low_T11Y69));
  sky130_fd_sc_hd__conb_1 conb_T11Y7 (.HI(tie_high_T11Y7), .LO(tie_low_T11Y7));
  sky130_fd_sc_hd__conb_1 conb_T11Y70 (.HI(tie_high_T11Y70), .LO(tie_low_T11Y70));
  sky130_fd_sc_hd__conb_1 conb_T11Y71 (.HI(tie_high_T11Y71), .LO(tie_low_T11Y71));
  sky130_fd_sc_hd__conb_1 conb_T11Y72 (.HI(tie_high_T11Y72), .LO(tie_low_T11Y72));
  sky130_fd_sc_hd__conb_1 conb_T11Y73 (.HI(tie_high_T11Y73), .LO(tie_low_T11Y73));
  sky130_fd_sc_hd__conb_1 conb_T11Y74 (.HI(tie_high_T11Y74), .LO(tie_low_T11Y74));
  sky130_fd_sc_hd__conb_1 conb_T11Y75 (.HI(tie_high_T11Y75), .LO(tie_low_T11Y75));
  sky130_fd_sc_hd__conb_1 conb_T11Y76 (.HI(tie_high_T11Y76), .LO(tie_low_T11Y76));
  sky130_fd_sc_hd__conb_1 conb_T11Y77 (.HI(tie_high_T11Y77), .LO(tie_low_T11Y77));
  sky130_fd_sc_hd__conb_1 conb_T11Y78 (.HI(tie_high_T11Y78), .LO(tie_low_T11Y78));
  sky130_fd_sc_hd__conb_1 conb_T11Y79 (.HI(tie_high_T11Y79), .LO(tie_low_T11Y79));
  sky130_fd_sc_hd__conb_1 conb_T11Y8 (.HI(tie_high_T11Y8), .LO(tie_low_T11Y8));
  sky130_fd_sc_hd__conb_1 conb_T11Y80 (.HI(tie_high_T11Y80), .LO(tie_low_T11Y80));
  sky130_fd_sc_hd__conb_1 conb_T11Y81 (.HI(tie_high_T11Y81), .LO(tie_low_T11Y81));
  sky130_fd_sc_hd__conb_1 conb_T11Y82 (.HI(tie_high_T11Y82), .LO(tie_low_T11Y82));
  sky130_fd_sc_hd__conb_1 conb_T11Y83 (.HI(tie_high_T11Y83), .LO(tie_low_T11Y83));
  sky130_fd_sc_hd__conb_1 conb_T11Y84 (.HI(tie_high_T11Y84), .LO(tie_low_T11Y84));
  sky130_fd_sc_hd__conb_1 conb_T11Y85 (.HI(tie_high_T11Y85), .LO(tie_low_T11Y85));
  sky130_fd_sc_hd__conb_1 conb_T11Y86 (.HI(tie_high_T11Y86), .LO(tie_low_T11Y86));
  sky130_fd_sc_hd__conb_1 conb_T11Y87 (.HI(tie_high_T11Y87), .LO(tie_low_T11Y87));
  sky130_fd_sc_hd__conb_1 conb_T11Y88 (.HI(tie_high_T11Y88), .LO(tie_low_T11Y88));
  sky130_fd_sc_hd__conb_1 conb_T11Y89 (.HI(tie_high_T11Y89), .LO(tie_low_T11Y89));
  sky130_fd_sc_hd__conb_1 conb_T11Y9 (.HI(tie_high_T11Y9), .LO(tie_low_T11Y9));
  sky130_fd_sc_hd__conb_1 conb_T12Y0 (.HI(tie_high_T12Y0), .LO(tie_low_T12Y0));
  sky130_fd_sc_hd__conb_1 conb_T12Y1 (.HI(tie_high_T12Y1), .LO(tie_low_T12Y1));
  sky130_fd_sc_hd__conb_1 conb_T12Y10 (.HI(tie_high_T12Y10), .LO(tie_low_T12Y10));
  sky130_fd_sc_hd__conb_1 conb_T12Y11 (.HI(tie_high_T12Y11), .LO(tie_low_T12Y11));
  sky130_fd_sc_hd__conb_1 conb_T12Y12 (.HI(tie_high_T12Y12), .LO(tie_low_T12Y12));
  sky130_fd_sc_hd__conb_1 conb_T12Y13 (.HI(tie_high_T12Y13), .LO(tie_low_T12Y13));
  sky130_fd_sc_hd__conb_1 conb_T12Y14 (.HI(tie_high_T12Y14), .LO(tie_low_T12Y14));
  sky130_fd_sc_hd__conb_1 conb_T12Y15 (.HI(tie_high_T12Y15), .LO(tie_low_T12Y15));
  sky130_fd_sc_hd__conb_1 conb_T12Y16 (.HI(tie_high_T12Y16), .LO(tie_low_T12Y16));
  sky130_fd_sc_hd__conb_1 conb_T12Y17 (.HI(tie_high_T12Y17), .LO(tie_low_T12Y17));
  sky130_fd_sc_hd__conb_1 conb_T12Y18 (.HI(tie_high_T12Y18), .LO(tie_low_T12Y18));
  sky130_fd_sc_hd__conb_1 conb_T12Y19 (.HI(tie_high_T12Y19), .LO(tie_low_T12Y19));
  sky130_fd_sc_hd__conb_1 conb_T12Y2 (.HI(tie_high_T12Y2), .LO(tie_low_T12Y2));
  sky130_fd_sc_hd__conb_1 conb_T12Y20 (.HI(tie_high_T12Y20), .LO(tie_low_T12Y20));
  sky130_fd_sc_hd__conb_1 conb_T12Y21 (.HI(tie_high_T12Y21), .LO(tie_low_T12Y21));
  sky130_fd_sc_hd__conb_1 conb_T12Y22 (.HI(tie_high_T12Y22), .LO(tie_low_T12Y22));
  sky130_fd_sc_hd__conb_1 conb_T12Y23 (.HI(tie_high_T12Y23), .LO(tie_low_T12Y23));
  sky130_fd_sc_hd__conb_1 conb_T12Y24 (.HI(tie_high_T12Y24), .LO(tie_low_T12Y24));
  sky130_fd_sc_hd__conb_1 conb_T12Y25 (.HI(tie_high_T12Y25), .LO(tie_low_T12Y25));
  sky130_fd_sc_hd__conb_1 conb_T12Y26 (.HI(tie_high_T12Y26), .LO(tie_low_T12Y26));
  sky130_fd_sc_hd__conb_1 conb_T12Y27 (.HI(tie_high_T12Y27), .LO(tie_low_T12Y27));
  sky130_fd_sc_hd__conb_1 conb_T12Y28 (.HI(tie_high_T12Y28), .LO(tie_low_T12Y28));
  sky130_fd_sc_hd__conb_1 conb_T12Y29 (.HI(tie_high_T12Y29), .LO(tie_low_T12Y29));
  sky130_fd_sc_hd__conb_1 conb_T12Y3 (.HI(tie_high_T12Y3), .LO(tie_low_T12Y3));
  sky130_fd_sc_hd__conb_1 conb_T12Y30 (.HI(tie_high_T12Y30), .LO(tie_low_T12Y30));
  sky130_fd_sc_hd__conb_1 conb_T12Y31 (.HI(tie_high_T12Y31), .LO(tie_low_T12Y31));
  sky130_fd_sc_hd__conb_1 conb_T12Y32 (.HI(tie_high_T12Y32), .LO(tie_low_T12Y32));
  sky130_fd_sc_hd__conb_1 conb_T12Y33 (.HI(tie_high_T12Y33), .LO(tie_low_T12Y33));
  sky130_fd_sc_hd__conb_1 conb_T12Y34 (.HI(tie_high_T12Y34), .LO(tie_low_T12Y34));
  sky130_fd_sc_hd__conb_1 conb_T12Y35 (.HI(tie_high_T12Y35), .LO(tie_low_T12Y35));
  sky130_fd_sc_hd__conb_1 conb_T12Y36 (.HI(tie_high_T12Y36), .LO(tie_low_T12Y36));
  sky130_fd_sc_hd__conb_1 conb_T12Y37 (.HI(tie_high_T12Y37), .LO(tie_low_T12Y37));
  sky130_fd_sc_hd__conb_1 conb_T12Y38 (.HI(tie_high_T12Y38), .LO(tie_low_T12Y38));
  sky130_fd_sc_hd__conb_1 conb_T12Y39 (.HI(tie_high_T12Y39), .LO(tie_low_T12Y39));
  sky130_fd_sc_hd__conb_1 conb_T12Y4 (.HI(tie_high_T12Y4), .LO(tie_low_T12Y4));
  sky130_fd_sc_hd__conb_1 conb_T12Y40 (.HI(tie_high_T12Y40), .LO(tie_low_T12Y40));
  sky130_fd_sc_hd__conb_1 conb_T12Y41 (.HI(tie_high_T12Y41), .LO(tie_low_T12Y41));
  sky130_fd_sc_hd__conb_1 conb_T12Y42 (.HI(tie_high_T12Y42), .LO(tie_low_T12Y42));
  sky130_fd_sc_hd__conb_1 conb_T12Y43 (.HI(tie_high_T12Y43), .LO(tie_low_T12Y43));
  sky130_fd_sc_hd__conb_1 conb_T12Y44 (.HI(tie_high_T12Y44), .LO(tie_low_T12Y44));
  sky130_fd_sc_hd__conb_1 conb_T12Y45 (.HI(tie_high_T12Y45), .LO(tie_low_T12Y45));
  sky130_fd_sc_hd__conb_1 conb_T12Y46 (.HI(tie_high_T12Y46), .LO(tie_low_T12Y46));
  sky130_fd_sc_hd__conb_1 conb_T12Y47 (.HI(tie_high_T12Y47), .LO(tie_low_T12Y47));
  sky130_fd_sc_hd__conb_1 conb_T12Y48 (.HI(tie_high_T12Y48), .LO(tie_low_T12Y48));
  sky130_fd_sc_hd__conb_1 conb_T12Y49 (.HI(tie_high_T12Y49), .LO(tie_low_T12Y49));
  sky130_fd_sc_hd__conb_1 conb_T12Y5 (.HI(tie_high_T12Y5), .LO(tie_low_T12Y5));
  sky130_fd_sc_hd__conb_1 conb_T12Y50 (.HI(tie_high_T12Y50), .LO(tie_low_T12Y50));
  sky130_fd_sc_hd__conb_1 conb_T12Y51 (.HI(tie_high_T12Y51), .LO(tie_low_T12Y51));
  sky130_fd_sc_hd__conb_1 conb_T12Y52 (.HI(tie_high_T12Y52), .LO(tie_low_T12Y52));
  sky130_fd_sc_hd__conb_1 conb_T12Y53 (.HI(tie_high_T12Y53), .LO(tie_low_T12Y53));
  sky130_fd_sc_hd__conb_1 conb_T12Y54 (.HI(tie_high_T12Y54), .LO(tie_low_T12Y54));
  sky130_fd_sc_hd__conb_1 conb_T12Y55 (.HI(tie_high_T12Y55), .LO(tie_low_T12Y55));
  sky130_fd_sc_hd__conb_1 conb_T12Y56 (.HI(tie_high_T12Y56), .LO(tie_low_T12Y56));
  sky130_fd_sc_hd__conb_1 conb_T12Y57 (.HI(tie_high_T12Y57), .LO(tie_low_T12Y57));
  sky130_fd_sc_hd__conb_1 conb_T12Y58 (.HI(tie_high_T12Y58), .LO(tie_low_T12Y58));
  sky130_fd_sc_hd__conb_1 conb_T12Y59 (.HI(tie_high_T12Y59), .LO(tie_low_T12Y59));
  sky130_fd_sc_hd__conb_1 conb_T12Y6 (.HI(tie_high_T12Y6), .LO(tie_low_T12Y6));
  sky130_fd_sc_hd__conb_1 conb_T12Y60 (.HI(tie_high_T12Y60), .LO(tie_low_T12Y60));
  sky130_fd_sc_hd__conb_1 conb_T12Y61 (.HI(tie_high_T12Y61), .LO(tie_low_T12Y61));
  sky130_fd_sc_hd__conb_1 conb_T12Y62 (.HI(tie_high_T12Y62), .LO(tie_low_T12Y62));
  sky130_fd_sc_hd__conb_1 conb_T12Y63 (.HI(tie_high_T12Y63), .LO(tie_low_T12Y63));
  sky130_fd_sc_hd__conb_1 conb_T12Y64 (.HI(tie_high_T12Y64), .LO(tie_low_T12Y64));
  sky130_fd_sc_hd__conb_1 conb_T12Y65 (.HI(tie_high_T12Y65), .LO(tie_low_T12Y65));
  sky130_fd_sc_hd__conb_1 conb_T12Y66 (.HI(tie_high_T12Y66), .LO(tie_low_T12Y66));
  sky130_fd_sc_hd__conb_1 conb_T12Y67 (.HI(tie_high_T12Y67), .LO(tie_low_T12Y67));
  sky130_fd_sc_hd__conb_1 conb_T12Y68 (.HI(tie_high_T12Y68), .LO(tie_low_T12Y68));
  sky130_fd_sc_hd__conb_1 conb_T12Y69 (.HI(tie_high_T12Y69), .LO(tie_low_T12Y69));
  sky130_fd_sc_hd__conb_1 conb_T12Y7 (.HI(tie_high_T12Y7), .LO(tie_low_T12Y7));
  sky130_fd_sc_hd__conb_1 conb_T12Y70 (.HI(tie_high_T12Y70), .LO(tie_low_T12Y70));
  sky130_fd_sc_hd__conb_1 conb_T12Y71 (.HI(tie_high_T12Y71), .LO(tie_low_T12Y71));
  sky130_fd_sc_hd__conb_1 conb_T12Y72 (.HI(tie_high_T12Y72), .LO(tie_low_T12Y72));
  sky130_fd_sc_hd__conb_1 conb_T12Y73 (.HI(tie_high_T12Y73), .LO(tie_low_T12Y73));
  sky130_fd_sc_hd__conb_1 conb_T12Y74 (.HI(tie_high_T12Y74), .LO(tie_low_T12Y74));
  sky130_fd_sc_hd__conb_1 conb_T12Y75 (.HI(tie_high_T12Y75), .LO(tie_low_T12Y75));
  sky130_fd_sc_hd__conb_1 conb_T12Y76 (.HI(tie_high_T12Y76), .LO(tie_low_T12Y76));
  sky130_fd_sc_hd__conb_1 conb_T12Y77 (.HI(tie_high_T12Y77), .LO(tie_low_T12Y77));
  sky130_fd_sc_hd__conb_1 conb_T12Y78 (.HI(tie_high_T12Y78), .LO(tie_low_T12Y78));
  sky130_fd_sc_hd__conb_1 conb_T12Y79 (.HI(tie_high_T12Y79), .LO(tie_low_T12Y79));
  sky130_fd_sc_hd__conb_1 conb_T12Y8 (.HI(tie_high_T12Y8), .LO(tie_low_T12Y8));
  sky130_fd_sc_hd__conb_1 conb_T12Y80 (.HI(tie_high_T12Y80), .LO(tie_low_T12Y80));
  sky130_fd_sc_hd__conb_1 conb_T12Y81 (.HI(tie_high_T12Y81), .LO(tie_low_T12Y81));
  sky130_fd_sc_hd__conb_1 conb_T12Y82 (.HI(tie_high_T12Y82), .LO(tie_low_T12Y82));
  sky130_fd_sc_hd__conb_1 conb_T12Y83 (.HI(tie_high_T12Y83), .LO(tie_low_T12Y83));
  sky130_fd_sc_hd__conb_1 conb_T12Y84 (.HI(tie_high_T12Y84), .LO(tie_low_T12Y84));
  sky130_fd_sc_hd__conb_1 conb_T12Y85 (.HI(tie_high_T12Y85), .LO(tie_low_T12Y85));
  sky130_fd_sc_hd__conb_1 conb_T12Y86 (.HI(tie_high_T12Y86), .LO(tie_low_T12Y86));
  sky130_fd_sc_hd__conb_1 conb_T12Y87 (.HI(tie_high_T12Y87), .LO(tie_low_T12Y87));
  sky130_fd_sc_hd__conb_1 conb_T12Y88 (.HI(tie_high_T12Y88), .LO(tie_low_T12Y88));
  sky130_fd_sc_hd__conb_1 conb_T12Y89 (.HI(tie_high_T12Y89), .LO(tie_low_T12Y89));
  sky130_fd_sc_hd__conb_1 conb_T12Y9 (.HI(tie_high_T12Y9), .LO(tie_low_T12Y9));
  sky130_fd_sc_hd__conb_1 conb_T13Y0 (.HI(tie_high_T13Y0), .LO(tie_low_T13Y0));
  sky130_fd_sc_hd__conb_1 conb_T13Y1 (.HI(tie_high_T13Y1), .LO(tie_low_T13Y1));
  sky130_fd_sc_hd__conb_1 conb_T13Y10 (.HI(tie_high_T13Y10), .LO(tie_low_T13Y10));
  sky130_fd_sc_hd__conb_1 conb_T13Y11 (.HI(tie_high_T13Y11), .LO(tie_low_T13Y11));
  sky130_fd_sc_hd__conb_1 conb_T13Y12 (.HI(tie_high_T13Y12), .LO(tie_low_T13Y12));
  sky130_fd_sc_hd__conb_1 conb_T13Y13 (.HI(tie_high_T13Y13), .LO(tie_low_T13Y13));
  sky130_fd_sc_hd__conb_1 conb_T13Y14 (.HI(tie_high_T13Y14), .LO(tie_low_T13Y14));
  sky130_fd_sc_hd__conb_1 conb_T13Y15 (.HI(tie_high_T13Y15), .LO(tie_low_T13Y15));
  sky130_fd_sc_hd__conb_1 conb_T13Y16 (.HI(tie_high_T13Y16), .LO(tie_low_T13Y16));
  sky130_fd_sc_hd__conb_1 conb_T13Y17 (.HI(tie_high_T13Y17), .LO(tie_low_T13Y17));
  sky130_fd_sc_hd__conb_1 conb_T13Y18 (.HI(tie_high_T13Y18), .LO(tie_low_T13Y18));
  sky130_fd_sc_hd__conb_1 conb_T13Y19 (.HI(tie_high_T13Y19), .LO(tie_low_T13Y19));
  sky130_fd_sc_hd__conb_1 conb_T13Y2 (.HI(tie_high_T13Y2), .LO(tie_low_T13Y2));
  sky130_fd_sc_hd__conb_1 conb_T13Y20 (.HI(tie_high_T13Y20), .LO(tie_low_T13Y20));
  sky130_fd_sc_hd__conb_1 conb_T13Y21 (.HI(tie_high_T13Y21), .LO(tie_low_T13Y21));
  sky130_fd_sc_hd__conb_1 conb_T13Y22 (.HI(tie_high_T13Y22), .LO(tie_low_T13Y22));
  sky130_fd_sc_hd__conb_1 conb_T13Y23 (.HI(tie_high_T13Y23), .LO(tie_low_T13Y23));
  sky130_fd_sc_hd__conb_1 conb_T13Y24 (.HI(tie_high_T13Y24), .LO(tie_low_T13Y24));
  sky130_fd_sc_hd__conb_1 conb_T13Y25 (.HI(tie_high_T13Y25), .LO(tie_low_T13Y25));
  sky130_fd_sc_hd__conb_1 conb_T13Y26 (.HI(tie_high_T13Y26), .LO(tie_low_T13Y26));
  sky130_fd_sc_hd__conb_1 conb_T13Y27 (.HI(tie_high_T13Y27), .LO(tie_low_T13Y27));
  sky130_fd_sc_hd__conb_1 conb_T13Y28 (.HI(tie_high_T13Y28), .LO(tie_low_T13Y28));
  sky130_fd_sc_hd__conb_1 conb_T13Y29 (.HI(tie_high_T13Y29), .LO(tie_low_T13Y29));
  sky130_fd_sc_hd__conb_1 conb_T13Y3 (.HI(tie_high_T13Y3), .LO(tie_low_T13Y3));
  sky130_fd_sc_hd__conb_1 conb_T13Y30 (.HI(tie_high_T13Y30), .LO(tie_low_T13Y30));
  sky130_fd_sc_hd__conb_1 conb_T13Y31 (.HI(tie_high_T13Y31), .LO(tie_low_T13Y31));
  sky130_fd_sc_hd__conb_1 conb_T13Y32 (.HI(tie_high_T13Y32), .LO(tie_low_T13Y32));
  sky130_fd_sc_hd__conb_1 conb_T13Y33 (.HI(tie_high_T13Y33), .LO(tie_low_T13Y33));
  sky130_fd_sc_hd__conb_1 conb_T13Y34 (.HI(tie_high_T13Y34), .LO(tie_low_T13Y34));
  sky130_fd_sc_hd__conb_1 conb_T13Y35 (.HI(tie_high_T13Y35), .LO(tie_low_T13Y35));
  sky130_fd_sc_hd__conb_1 conb_T13Y36 (.HI(tie_high_T13Y36), .LO(tie_low_T13Y36));
  sky130_fd_sc_hd__conb_1 conb_T13Y37 (.HI(tie_high_T13Y37), .LO(tie_low_T13Y37));
  sky130_fd_sc_hd__conb_1 conb_T13Y38 (.HI(tie_high_T13Y38), .LO(tie_low_T13Y38));
  sky130_fd_sc_hd__conb_1 conb_T13Y39 (.HI(tie_high_T13Y39), .LO(tie_low_T13Y39));
  sky130_fd_sc_hd__conb_1 conb_T13Y4 (.HI(tie_high_T13Y4), .LO(tie_low_T13Y4));
  sky130_fd_sc_hd__conb_1 conb_T13Y40 (.HI(tie_high_T13Y40), .LO(tie_low_T13Y40));
  sky130_fd_sc_hd__conb_1 conb_T13Y41 (.HI(tie_high_T13Y41), .LO(tie_low_T13Y41));
  sky130_fd_sc_hd__conb_1 conb_T13Y42 (.HI(tie_high_T13Y42), .LO(tie_low_T13Y42));
  sky130_fd_sc_hd__conb_1 conb_T13Y43 (.HI(tie_high_T13Y43), .LO(tie_low_T13Y43));
  sky130_fd_sc_hd__conb_1 conb_T13Y44 (.HI(tie_high_T13Y44), .LO(tie_low_T13Y44));
  sky130_fd_sc_hd__conb_1 conb_T13Y45 (.HI(tie_high_T13Y45), .LO(tie_low_T13Y45));
  sky130_fd_sc_hd__conb_1 conb_T13Y46 (.HI(tie_high_T13Y46), .LO(tie_low_T13Y46));
  sky130_fd_sc_hd__conb_1 conb_T13Y47 (.HI(tie_high_T13Y47), .LO(tie_low_T13Y47));
  sky130_fd_sc_hd__conb_1 conb_T13Y48 (.HI(tie_high_T13Y48), .LO(tie_low_T13Y48));
  sky130_fd_sc_hd__conb_1 conb_T13Y49 (.HI(tie_high_T13Y49), .LO(tie_low_T13Y49));
  sky130_fd_sc_hd__conb_1 conb_T13Y5 (.HI(tie_high_T13Y5), .LO(tie_low_T13Y5));
  sky130_fd_sc_hd__conb_1 conb_T13Y50 (.HI(tie_high_T13Y50), .LO(tie_low_T13Y50));
  sky130_fd_sc_hd__conb_1 conb_T13Y51 (.HI(tie_high_T13Y51), .LO(tie_low_T13Y51));
  sky130_fd_sc_hd__conb_1 conb_T13Y52 (.HI(tie_high_T13Y52), .LO(tie_low_T13Y52));
  sky130_fd_sc_hd__conb_1 conb_T13Y53 (.HI(tie_high_T13Y53), .LO(tie_low_T13Y53));
  sky130_fd_sc_hd__conb_1 conb_T13Y54 (.HI(tie_high_T13Y54), .LO(tie_low_T13Y54));
  sky130_fd_sc_hd__conb_1 conb_T13Y55 (.HI(tie_high_T13Y55), .LO(tie_low_T13Y55));
  sky130_fd_sc_hd__conb_1 conb_T13Y56 (.HI(tie_high_T13Y56), .LO(tie_low_T13Y56));
  sky130_fd_sc_hd__conb_1 conb_T13Y57 (.HI(tie_high_T13Y57), .LO(tie_low_T13Y57));
  sky130_fd_sc_hd__conb_1 conb_T13Y58 (.HI(tie_high_T13Y58), .LO(tie_low_T13Y58));
  sky130_fd_sc_hd__conb_1 conb_T13Y59 (.HI(tie_high_T13Y59), .LO(tie_low_T13Y59));
  sky130_fd_sc_hd__conb_1 conb_T13Y6 (.HI(tie_high_T13Y6), .LO(tie_low_T13Y6));
  sky130_fd_sc_hd__conb_1 conb_T13Y60 (.HI(tie_high_T13Y60), .LO(tie_low_T13Y60));
  sky130_fd_sc_hd__conb_1 conb_T13Y61 (.HI(tie_high_T13Y61), .LO(tie_low_T13Y61));
  sky130_fd_sc_hd__conb_1 conb_T13Y62 (.HI(tie_high_T13Y62), .LO(tie_low_T13Y62));
  sky130_fd_sc_hd__conb_1 conb_T13Y63 (.HI(tie_high_T13Y63), .LO(tie_low_T13Y63));
  sky130_fd_sc_hd__conb_1 conb_T13Y64 (.HI(tie_high_T13Y64), .LO(tie_low_T13Y64));
  sky130_fd_sc_hd__conb_1 conb_T13Y65 (.HI(tie_high_T13Y65), .LO(tie_low_T13Y65));
  sky130_fd_sc_hd__conb_1 conb_T13Y66 (.HI(tie_high_T13Y66), .LO(tie_low_T13Y66));
  sky130_fd_sc_hd__conb_1 conb_T13Y67 (.HI(tie_high_T13Y67), .LO(tie_low_T13Y67));
  sky130_fd_sc_hd__conb_1 conb_T13Y68 (.HI(tie_high_T13Y68), .LO(tie_low_T13Y68));
  sky130_fd_sc_hd__conb_1 conb_T13Y69 (.HI(tie_high_T13Y69), .LO(tie_low_T13Y69));
  sky130_fd_sc_hd__conb_1 conb_T13Y7 (.HI(tie_high_T13Y7), .LO(tie_low_T13Y7));
  sky130_fd_sc_hd__conb_1 conb_T13Y70 (.HI(tie_high_T13Y70), .LO(tie_low_T13Y70));
  sky130_fd_sc_hd__conb_1 conb_T13Y71 (.HI(tie_high_T13Y71), .LO(tie_low_T13Y71));
  sky130_fd_sc_hd__conb_1 conb_T13Y72 (.HI(tie_high_T13Y72), .LO(tie_low_T13Y72));
  sky130_fd_sc_hd__conb_1 conb_T13Y73 (.HI(tie_high_T13Y73), .LO(tie_low_T13Y73));
  sky130_fd_sc_hd__conb_1 conb_T13Y74 (.HI(tie_high_T13Y74), .LO(tie_low_T13Y74));
  sky130_fd_sc_hd__conb_1 conb_T13Y75 (.HI(tie_high_T13Y75), .LO(tie_low_T13Y75));
  sky130_fd_sc_hd__conb_1 conb_T13Y76 (.HI(tie_high_T13Y76), .LO(tie_low_T13Y76));
  sky130_fd_sc_hd__conb_1 conb_T13Y77 (.HI(tie_high_T13Y77), .LO(tie_low_T13Y77));
  sky130_fd_sc_hd__conb_1 conb_T13Y78 (.HI(tie_high_T13Y78), .LO(tie_low_T13Y78));
  sky130_fd_sc_hd__conb_1 conb_T13Y79 (.HI(tie_high_T13Y79), .LO(tie_low_T13Y79));
  sky130_fd_sc_hd__conb_1 conb_T13Y8 (.HI(tie_high_T13Y8), .LO(tie_low_T13Y8));
  sky130_fd_sc_hd__conb_1 conb_T13Y80 (.HI(tie_high_T13Y80), .LO(tie_low_T13Y80));
  sky130_fd_sc_hd__conb_1 conb_T13Y81 (.HI(tie_high_T13Y81), .LO(tie_low_T13Y81));
  sky130_fd_sc_hd__conb_1 conb_T13Y82 (.HI(tie_high_T13Y82), .LO(tie_low_T13Y82));
  sky130_fd_sc_hd__conb_1 conb_T13Y83 (.HI(tie_high_T13Y83), .LO(tie_low_T13Y83));
  sky130_fd_sc_hd__conb_1 conb_T13Y84 (.HI(tie_high_T13Y84), .LO(tie_low_T13Y84));
  sky130_fd_sc_hd__conb_1 conb_T13Y85 (.HI(tie_high_T13Y85), .LO(tie_low_T13Y85));
  sky130_fd_sc_hd__conb_1 conb_T13Y86 (.HI(tie_high_T13Y86), .LO(tie_low_T13Y86));
  sky130_fd_sc_hd__conb_1 conb_T13Y87 (.HI(tie_high_T13Y87), .LO(tie_low_T13Y87));
  sky130_fd_sc_hd__conb_1 conb_T13Y88 (.HI(tie_high_T13Y88), .LO(tie_low_T13Y88));
  sky130_fd_sc_hd__conb_1 conb_T13Y89 (.HI(tie_high_T13Y89), .LO(tie_low_T13Y89));
  sky130_fd_sc_hd__conb_1 conb_T13Y9 (.HI(tie_high_T13Y9), .LO(tie_low_T13Y9));
  sky130_fd_sc_hd__conb_1 conb_T14Y0 (.HI(tie_high_T14Y0), .LO(tie_low_T14Y0));
  sky130_fd_sc_hd__conb_1 conb_T14Y1 (.HI(tie_high_T14Y1), .LO(tie_low_T14Y1));
  sky130_fd_sc_hd__conb_1 conb_T14Y10 (.HI(tie_high_T14Y10), .LO(tie_low_T14Y10));
  sky130_fd_sc_hd__conb_1 conb_T14Y11 (.HI(tie_high_T14Y11), .LO(tie_low_T14Y11));
  sky130_fd_sc_hd__conb_1 conb_T14Y12 (.HI(tie_high_T14Y12), .LO(tie_low_T14Y12));
  sky130_fd_sc_hd__conb_1 conb_T14Y13 (.HI(tie_high_T14Y13), .LO(tie_low_T14Y13));
  sky130_fd_sc_hd__conb_1 conb_T14Y14 (.HI(tie_high_T14Y14), .LO(tie_low_T14Y14));
  sky130_fd_sc_hd__conb_1 conb_T14Y15 (.HI(tie_high_T14Y15), .LO(tie_low_T14Y15));
  sky130_fd_sc_hd__conb_1 conb_T14Y16 (.HI(tie_high_T14Y16), .LO(tie_low_T14Y16));
  sky130_fd_sc_hd__conb_1 conb_T14Y17 (.HI(tie_high_T14Y17), .LO(tie_low_T14Y17));
  sky130_fd_sc_hd__conb_1 conb_T14Y18 (.HI(tie_high_T14Y18), .LO(tie_low_T14Y18));
  sky130_fd_sc_hd__conb_1 conb_T14Y19 (.HI(tie_high_T14Y19), .LO(tie_low_T14Y19));
  sky130_fd_sc_hd__conb_1 conb_T14Y2 (.HI(tie_high_T14Y2), .LO(tie_low_T14Y2));
  sky130_fd_sc_hd__conb_1 conb_T14Y20 (.HI(tie_high_T14Y20), .LO(tie_low_T14Y20));
  sky130_fd_sc_hd__conb_1 conb_T14Y21 (.HI(tie_high_T14Y21), .LO(tie_low_T14Y21));
  sky130_fd_sc_hd__conb_1 conb_T14Y22 (.HI(tie_high_T14Y22), .LO(tie_low_T14Y22));
  sky130_fd_sc_hd__conb_1 conb_T14Y23 (.HI(tie_high_T14Y23), .LO(tie_low_T14Y23));
  sky130_fd_sc_hd__conb_1 conb_T14Y24 (.HI(tie_high_T14Y24), .LO(tie_low_T14Y24));
  sky130_fd_sc_hd__conb_1 conb_T14Y25 (.HI(tie_high_T14Y25), .LO(tie_low_T14Y25));
  sky130_fd_sc_hd__conb_1 conb_T14Y26 (.HI(tie_high_T14Y26), .LO(tie_low_T14Y26));
  sky130_fd_sc_hd__conb_1 conb_T14Y27 (.HI(tie_high_T14Y27), .LO(tie_low_T14Y27));
  sky130_fd_sc_hd__conb_1 conb_T14Y28 (.HI(tie_high_T14Y28), .LO(tie_low_T14Y28));
  sky130_fd_sc_hd__conb_1 conb_T14Y29 (.HI(tie_high_T14Y29), .LO(tie_low_T14Y29));
  sky130_fd_sc_hd__conb_1 conb_T14Y3 (.HI(tie_high_T14Y3), .LO(tie_low_T14Y3));
  sky130_fd_sc_hd__conb_1 conb_T14Y30 (.HI(tie_high_T14Y30), .LO(tie_low_T14Y30));
  sky130_fd_sc_hd__conb_1 conb_T14Y31 (.HI(tie_high_T14Y31), .LO(tie_low_T14Y31));
  sky130_fd_sc_hd__conb_1 conb_T14Y32 (.HI(tie_high_T14Y32), .LO(tie_low_T14Y32));
  sky130_fd_sc_hd__conb_1 conb_T14Y33 (.HI(tie_high_T14Y33), .LO(tie_low_T14Y33));
  sky130_fd_sc_hd__conb_1 conb_T14Y34 (.HI(tie_high_T14Y34), .LO(tie_low_T14Y34));
  sky130_fd_sc_hd__conb_1 conb_T14Y35 (.HI(tie_high_T14Y35), .LO(tie_low_T14Y35));
  sky130_fd_sc_hd__conb_1 conb_T14Y36 (.HI(tie_high_T14Y36), .LO(tie_low_T14Y36));
  sky130_fd_sc_hd__conb_1 conb_T14Y37 (.HI(tie_high_T14Y37), .LO(tie_low_T14Y37));
  sky130_fd_sc_hd__conb_1 conb_T14Y38 (.HI(tie_high_T14Y38), .LO(tie_low_T14Y38));
  sky130_fd_sc_hd__conb_1 conb_T14Y39 (.HI(tie_high_T14Y39), .LO(tie_low_T14Y39));
  sky130_fd_sc_hd__conb_1 conb_T14Y4 (.HI(tie_high_T14Y4), .LO(tie_low_T14Y4));
  sky130_fd_sc_hd__conb_1 conb_T14Y40 (.HI(tie_high_T14Y40), .LO(tie_low_T14Y40));
  sky130_fd_sc_hd__conb_1 conb_T14Y41 (.HI(tie_high_T14Y41), .LO(tie_low_T14Y41));
  sky130_fd_sc_hd__conb_1 conb_T14Y42 (.HI(tie_high_T14Y42), .LO(tie_low_T14Y42));
  sky130_fd_sc_hd__conb_1 conb_T14Y43 (.HI(tie_high_T14Y43), .LO(tie_low_T14Y43));
  sky130_fd_sc_hd__conb_1 conb_T14Y44 (.HI(tie_high_T14Y44), .LO(tie_low_T14Y44));
  sky130_fd_sc_hd__conb_1 conb_T14Y45 (.HI(tie_high_T14Y45), .LO(tie_low_T14Y45));
  sky130_fd_sc_hd__conb_1 conb_T14Y46 (.HI(tie_high_T14Y46), .LO(tie_low_T14Y46));
  sky130_fd_sc_hd__conb_1 conb_T14Y47 (.HI(tie_high_T14Y47), .LO(tie_low_T14Y47));
  sky130_fd_sc_hd__conb_1 conb_T14Y48 (.HI(tie_high_T14Y48), .LO(tie_low_T14Y48));
  sky130_fd_sc_hd__conb_1 conb_T14Y49 (.HI(tie_high_T14Y49), .LO(tie_low_T14Y49));
  sky130_fd_sc_hd__conb_1 conb_T14Y5 (.HI(tie_high_T14Y5), .LO(tie_low_T14Y5));
  sky130_fd_sc_hd__conb_1 conb_T14Y50 (.HI(tie_high_T14Y50), .LO(tie_low_T14Y50));
  sky130_fd_sc_hd__conb_1 conb_T14Y51 (.HI(tie_high_T14Y51), .LO(tie_low_T14Y51));
  sky130_fd_sc_hd__conb_1 conb_T14Y52 (.HI(tie_high_T14Y52), .LO(tie_low_T14Y52));
  sky130_fd_sc_hd__conb_1 conb_T14Y53 (.HI(tie_high_T14Y53), .LO(tie_low_T14Y53));
  sky130_fd_sc_hd__conb_1 conb_T14Y54 (.HI(tie_high_T14Y54), .LO(tie_low_T14Y54));
  sky130_fd_sc_hd__conb_1 conb_T14Y55 (.HI(tie_high_T14Y55), .LO(tie_low_T14Y55));
  sky130_fd_sc_hd__conb_1 conb_T14Y56 (.HI(tie_high_T14Y56), .LO(tie_low_T14Y56));
  sky130_fd_sc_hd__conb_1 conb_T14Y57 (.HI(tie_high_T14Y57), .LO(tie_low_T14Y57));
  sky130_fd_sc_hd__conb_1 conb_T14Y58 (.HI(tie_high_T14Y58), .LO(tie_low_T14Y58));
  sky130_fd_sc_hd__conb_1 conb_T14Y59 (.HI(tie_high_T14Y59), .LO(tie_low_T14Y59));
  sky130_fd_sc_hd__conb_1 conb_T14Y6 (.HI(tie_high_T14Y6), .LO(tie_low_T14Y6));
  sky130_fd_sc_hd__conb_1 conb_T14Y60 (.HI(tie_high_T14Y60), .LO(tie_low_T14Y60));
  sky130_fd_sc_hd__conb_1 conb_T14Y61 (.HI(tie_high_T14Y61), .LO(tie_low_T14Y61));
  sky130_fd_sc_hd__conb_1 conb_T14Y62 (.HI(tie_high_T14Y62), .LO(tie_low_T14Y62));
  sky130_fd_sc_hd__conb_1 conb_T14Y63 (.HI(tie_high_T14Y63), .LO(tie_low_T14Y63));
  sky130_fd_sc_hd__conb_1 conb_T14Y64 (.HI(tie_high_T14Y64), .LO(tie_low_T14Y64));
  sky130_fd_sc_hd__conb_1 conb_T14Y65 (.HI(tie_high_T14Y65), .LO(tie_low_T14Y65));
  sky130_fd_sc_hd__conb_1 conb_T14Y66 (.HI(tie_high_T14Y66), .LO(tie_low_T14Y66));
  sky130_fd_sc_hd__conb_1 conb_T14Y67 (.HI(tie_high_T14Y67), .LO(tie_low_T14Y67));
  sky130_fd_sc_hd__conb_1 conb_T14Y68 (.HI(tie_high_T14Y68), .LO(tie_low_T14Y68));
  sky130_fd_sc_hd__conb_1 conb_T14Y69 (.HI(tie_high_T14Y69), .LO(tie_low_T14Y69));
  sky130_fd_sc_hd__conb_1 conb_T14Y7 (.HI(tie_high_T14Y7), .LO(tie_low_T14Y7));
  sky130_fd_sc_hd__conb_1 conb_T14Y70 (.HI(tie_high_T14Y70), .LO(tie_low_T14Y70));
  sky130_fd_sc_hd__conb_1 conb_T14Y71 (.HI(tie_high_T14Y71), .LO(tie_low_T14Y71));
  sky130_fd_sc_hd__conb_1 conb_T14Y72 (.HI(tie_high_T14Y72), .LO(tie_low_T14Y72));
  sky130_fd_sc_hd__conb_1 conb_T14Y73 (.HI(tie_high_T14Y73), .LO(tie_low_T14Y73));
  sky130_fd_sc_hd__conb_1 conb_T14Y74 (.HI(tie_high_T14Y74), .LO(tie_low_T14Y74));
  sky130_fd_sc_hd__conb_1 conb_T14Y75 (.HI(tie_high_T14Y75), .LO(tie_low_T14Y75));
  sky130_fd_sc_hd__conb_1 conb_T14Y76 (.HI(tie_high_T14Y76), .LO(tie_low_T14Y76));
  sky130_fd_sc_hd__conb_1 conb_T14Y77 (.HI(tie_high_T14Y77), .LO(tie_low_T14Y77));
  sky130_fd_sc_hd__conb_1 conb_T14Y78 (.HI(tie_high_T14Y78), .LO(tie_low_T14Y78));
  sky130_fd_sc_hd__conb_1 conb_T14Y79 (.HI(tie_high_T14Y79), .LO(tie_low_T14Y79));
  sky130_fd_sc_hd__conb_1 conb_T14Y8 (.HI(tie_high_T14Y8), .LO(tie_low_T14Y8));
  sky130_fd_sc_hd__conb_1 conb_T14Y80 (.HI(tie_high_T14Y80), .LO(tie_low_T14Y80));
  sky130_fd_sc_hd__conb_1 conb_T14Y81 (.HI(tie_high_T14Y81), .LO(tie_low_T14Y81));
  sky130_fd_sc_hd__conb_1 conb_T14Y82 (.HI(tie_high_T14Y82), .LO(tie_low_T14Y82));
  sky130_fd_sc_hd__conb_1 conb_T14Y83 (.HI(tie_high_T14Y83), .LO(tie_low_T14Y83));
  sky130_fd_sc_hd__conb_1 conb_T14Y84 (.HI(tie_high_T14Y84), .LO(tie_low_T14Y84));
  sky130_fd_sc_hd__conb_1 conb_T14Y85 (.HI(tie_high_T14Y85), .LO(tie_low_T14Y85));
  sky130_fd_sc_hd__conb_1 conb_T14Y86 (.HI(tie_high_T14Y86), .LO(tie_low_T14Y86));
  sky130_fd_sc_hd__conb_1 conb_T14Y87 (.HI(tie_high_T14Y87), .LO(tie_low_T14Y87));
  sky130_fd_sc_hd__conb_1 conb_T14Y88 (.HI(tie_high_T14Y88), .LO(tie_low_T14Y88));
  sky130_fd_sc_hd__conb_1 conb_T14Y89 (.HI(tie_high_T14Y89), .LO(tie_low_T14Y89));
  sky130_fd_sc_hd__conb_1 conb_T14Y9 (.HI(tie_high_T14Y9), .LO(tie_low_T14Y9));
  sky130_fd_sc_hd__conb_1 conb_T15Y0 (.HI(tie_high_T15Y0), .LO(tie_low_T15Y0));
  sky130_fd_sc_hd__conb_1 conb_T15Y1 (.HI(tie_high_T15Y1), .LO(tie_low_T15Y1));
  sky130_fd_sc_hd__conb_1 conb_T15Y10 (.HI(tie_high_T15Y10), .LO(tie_low_T15Y10));
  sky130_fd_sc_hd__conb_1 conb_T15Y11 (.HI(tie_high_T15Y11), .LO(tie_low_T15Y11));
  sky130_fd_sc_hd__conb_1 conb_T15Y12 (.HI(tie_high_T15Y12), .LO(tie_low_T15Y12));
  sky130_fd_sc_hd__conb_1 conb_T15Y13 (.HI(tie_high_T15Y13), .LO(tie_low_T15Y13));
  sky130_fd_sc_hd__conb_1 conb_T15Y14 (.HI(tie_high_T15Y14), .LO(tie_low_T15Y14));
  sky130_fd_sc_hd__conb_1 conb_T15Y15 (.HI(tie_high_T15Y15), .LO(tie_low_T15Y15));
  sky130_fd_sc_hd__conb_1 conb_T15Y16 (.HI(tie_high_T15Y16), .LO(tie_low_T15Y16));
  sky130_fd_sc_hd__conb_1 conb_T15Y17 (.HI(tie_high_T15Y17), .LO(tie_low_T15Y17));
  sky130_fd_sc_hd__conb_1 conb_T15Y18 (.HI(tie_high_T15Y18), .LO(tie_low_T15Y18));
  sky130_fd_sc_hd__conb_1 conb_T15Y19 (.HI(tie_high_T15Y19), .LO(tie_low_T15Y19));
  sky130_fd_sc_hd__conb_1 conb_T15Y2 (.HI(tie_high_T15Y2), .LO(tie_low_T15Y2));
  sky130_fd_sc_hd__conb_1 conb_T15Y20 (.HI(tie_high_T15Y20), .LO(tie_low_T15Y20));
  sky130_fd_sc_hd__conb_1 conb_T15Y21 (.HI(tie_high_T15Y21), .LO(tie_low_T15Y21));
  sky130_fd_sc_hd__conb_1 conb_T15Y22 (.HI(tie_high_T15Y22), .LO(tie_low_T15Y22));
  sky130_fd_sc_hd__conb_1 conb_T15Y23 (.HI(tie_high_T15Y23), .LO(tie_low_T15Y23));
  sky130_fd_sc_hd__conb_1 conb_T15Y24 (.HI(tie_high_T15Y24), .LO(tie_low_T15Y24));
  sky130_fd_sc_hd__conb_1 conb_T15Y25 (.HI(tie_high_T15Y25), .LO(tie_low_T15Y25));
  sky130_fd_sc_hd__conb_1 conb_T15Y26 (.HI(tie_high_T15Y26), .LO(tie_low_T15Y26));
  sky130_fd_sc_hd__conb_1 conb_T15Y27 (.HI(tie_high_T15Y27), .LO(tie_low_T15Y27));
  sky130_fd_sc_hd__conb_1 conb_T15Y28 (.HI(tie_high_T15Y28), .LO(tie_low_T15Y28));
  sky130_fd_sc_hd__conb_1 conb_T15Y29 (.HI(tie_high_T15Y29), .LO(tie_low_T15Y29));
  sky130_fd_sc_hd__conb_1 conb_T15Y3 (.HI(tie_high_T15Y3), .LO(tie_low_T15Y3));
  sky130_fd_sc_hd__conb_1 conb_T15Y30 (.HI(tie_high_T15Y30), .LO(tie_low_T15Y30));
  sky130_fd_sc_hd__conb_1 conb_T15Y31 (.HI(tie_high_T15Y31), .LO(tie_low_T15Y31));
  sky130_fd_sc_hd__conb_1 conb_T15Y32 (.HI(tie_high_T15Y32), .LO(tie_low_T15Y32));
  sky130_fd_sc_hd__conb_1 conb_T15Y33 (.HI(tie_high_T15Y33), .LO(tie_low_T15Y33));
  sky130_fd_sc_hd__conb_1 conb_T15Y34 (.HI(tie_high_T15Y34), .LO(tie_low_T15Y34));
  sky130_fd_sc_hd__conb_1 conb_T15Y35 (.HI(tie_high_T15Y35), .LO(tie_low_T15Y35));
  sky130_fd_sc_hd__conb_1 conb_T15Y36 (.HI(tie_high_T15Y36), .LO(tie_low_T15Y36));
  sky130_fd_sc_hd__conb_1 conb_T15Y37 (.HI(tie_high_T15Y37), .LO(tie_low_T15Y37));
  sky130_fd_sc_hd__conb_1 conb_T15Y38 (.HI(tie_high_T15Y38), .LO(tie_low_T15Y38));
  sky130_fd_sc_hd__conb_1 conb_T15Y39 (.HI(tie_high_T15Y39), .LO(tie_low_T15Y39));
  sky130_fd_sc_hd__conb_1 conb_T15Y4 (.HI(tie_high_T15Y4), .LO(tie_low_T15Y4));
  sky130_fd_sc_hd__conb_1 conb_T15Y40 (.HI(tie_high_T15Y40), .LO(tie_low_T15Y40));
  sky130_fd_sc_hd__conb_1 conb_T15Y41 (.HI(tie_high_T15Y41), .LO(tie_low_T15Y41));
  sky130_fd_sc_hd__conb_1 conb_T15Y42 (.HI(tie_high_T15Y42), .LO(tie_low_T15Y42));
  sky130_fd_sc_hd__conb_1 conb_T15Y43 (.HI(tie_high_T15Y43), .LO(tie_low_T15Y43));
  sky130_fd_sc_hd__conb_1 conb_T15Y44 (.HI(tie_high_T15Y44), .LO(tie_low_T15Y44));
  sky130_fd_sc_hd__conb_1 conb_T15Y45 (.HI(tie_high_T15Y45), .LO(tie_low_T15Y45));
  sky130_fd_sc_hd__conb_1 conb_T15Y46 (.HI(tie_high_T15Y46), .LO(tie_low_T15Y46));
  sky130_fd_sc_hd__conb_1 conb_T15Y47 (.HI(tie_high_T15Y47), .LO(tie_low_T15Y47));
  sky130_fd_sc_hd__conb_1 conb_T15Y48 (.HI(tie_high_T15Y48), .LO(tie_low_T15Y48));
  sky130_fd_sc_hd__conb_1 conb_T15Y49 (.HI(tie_high_T15Y49), .LO(tie_low_T15Y49));
  sky130_fd_sc_hd__conb_1 conb_T15Y5 (.HI(tie_high_T15Y5), .LO(tie_low_T15Y5));
  sky130_fd_sc_hd__conb_1 conb_T15Y50 (.HI(tie_high_T15Y50), .LO(tie_low_T15Y50));
  sky130_fd_sc_hd__conb_1 conb_T15Y51 (.HI(tie_high_T15Y51), .LO(tie_low_T15Y51));
  sky130_fd_sc_hd__conb_1 conb_T15Y52 (.HI(tie_high_T15Y52), .LO(tie_low_T15Y52));
  sky130_fd_sc_hd__conb_1 conb_T15Y53 (.HI(tie_high_T15Y53), .LO(tie_low_T15Y53));
  sky130_fd_sc_hd__conb_1 conb_T15Y54 (.HI(tie_high_T15Y54), .LO(tie_low_T15Y54));
  sky130_fd_sc_hd__conb_1 conb_T15Y55 (.HI(tie_high_T15Y55), .LO(tie_low_T15Y55));
  sky130_fd_sc_hd__conb_1 conb_T15Y56 (.HI(tie_high_T15Y56), .LO(tie_low_T15Y56));
  sky130_fd_sc_hd__conb_1 conb_T15Y57 (.HI(tie_high_T15Y57), .LO(tie_low_T15Y57));
  sky130_fd_sc_hd__conb_1 conb_T15Y58 (.HI(tie_high_T15Y58), .LO(tie_low_T15Y58));
  sky130_fd_sc_hd__conb_1 conb_T15Y59 (.HI(tie_high_T15Y59), .LO(tie_low_T15Y59));
  sky130_fd_sc_hd__conb_1 conb_T15Y6 (.HI(tie_high_T15Y6), .LO(tie_low_T15Y6));
  sky130_fd_sc_hd__conb_1 conb_T15Y60 (.HI(tie_high_T15Y60), .LO(tie_low_T15Y60));
  sky130_fd_sc_hd__conb_1 conb_T15Y61 (.HI(tie_high_T15Y61), .LO(tie_low_T15Y61));
  sky130_fd_sc_hd__conb_1 conb_T15Y62 (.HI(tie_high_T15Y62), .LO(tie_low_T15Y62));
  sky130_fd_sc_hd__conb_1 conb_T15Y63 (.HI(tie_high_T15Y63), .LO(tie_low_T15Y63));
  sky130_fd_sc_hd__conb_1 conb_T15Y64 (.HI(tie_high_T15Y64), .LO(tie_low_T15Y64));
  sky130_fd_sc_hd__conb_1 conb_T15Y65 (.HI(tie_high_T15Y65), .LO(tie_low_T15Y65));
  sky130_fd_sc_hd__conb_1 conb_T15Y66 (.HI(tie_high_T15Y66), .LO(tie_low_T15Y66));
  sky130_fd_sc_hd__conb_1 conb_T15Y67 (.HI(tie_high_T15Y67), .LO(tie_low_T15Y67));
  sky130_fd_sc_hd__conb_1 conb_T15Y68 (.HI(tie_high_T15Y68), .LO(tie_low_T15Y68));
  sky130_fd_sc_hd__conb_1 conb_T15Y69 (.HI(tie_high_T15Y69), .LO(tie_low_T15Y69));
  sky130_fd_sc_hd__conb_1 conb_T15Y7 (.HI(tie_high_T15Y7), .LO(tie_low_T15Y7));
  sky130_fd_sc_hd__conb_1 conb_T15Y70 (.HI(tie_high_T15Y70), .LO(tie_low_T15Y70));
  sky130_fd_sc_hd__conb_1 conb_T15Y71 (.HI(tie_high_T15Y71), .LO(tie_low_T15Y71));
  sky130_fd_sc_hd__conb_1 conb_T15Y72 (.HI(tie_high_T15Y72), .LO(tie_low_T15Y72));
  sky130_fd_sc_hd__conb_1 conb_T15Y73 (.HI(tie_high_T15Y73), .LO(tie_low_T15Y73));
  sky130_fd_sc_hd__conb_1 conb_T15Y74 (.HI(tie_high_T15Y74), .LO(tie_low_T15Y74));
  sky130_fd_sc_hd__conb_1 conb_T15Y75 (.HI(tie_high_T15Y75), .LO(tie_low_T15Y75));
  sky130_fd_sc_hd__conb_1 conb_T15Y76 (.HI(tie_high_T15Y76), .LO(tie_low_T15Y76));
  sky130_fd_sc_hd__conb_1 conb_T15Y77 (.HI(tie_high_T15Y77), .LO(tie_low_T15Y77));
  sky130_fd_sc_hd__conb_1 conb_T15Y78 (.HI(tie_high_T15Y78), .LO(tie_low_T15Y78));
  sky130_fd_sc_hd__conb_1 conb_T15Y79 (.HI(tie_high_T15Y79), .LO(tie_low_T15Y79));
  sky130_fd_sc_hd__conb_1 conb_T15Y8 (.HI(tie_high_T15Y8), .LO(tie_low_T15Y8));
  sky130_fd_sc_hd__conb_1 conb_T15Y80 (.HI(tie_high_T15Y80), .LO(tie_low_T15Y80));
  sky130_fd_sc_hd__conb_1 conb_T15Y81 (.HI(tie_high_T15Y81), .LO(tie_low_T15Y81));
  sky130_fd_sc_hd__conb_1 conb_T15Y82 (.HI(tie_high_T15Y82), .LO(tie_low_T15Y82));
  sky130_fd_sc_hd__conb_1 conb_T15Y83 (.HI(tie_high_T15Y83), .LO(tie_low_T15Y83));
  sky130_fd_sc_hd__conb_1 conb_T15Y84 (.HI(tie_high_T15Y84), .LO(tie_low_T15Y84));
  sky130_fd_sc_hd__conb_1 conb_T15Y85 (.HI(tie_high_T15Y85), .LO(tie_low_T15Y85));
  sky130_fd_sc_hd__conb_1 conb_T15Y86 (.HI(tie_high_T15Y86), .LO(tie_low_T15Y86));
  sky130_fd_sc_hd__conb_1 conb_T15Y87 (.HI(tie_high_T15Y87), .LO(tie_low_T15Y87));
  sky130_fd_sc_hd__conb_1 conb_T15Y88 (.HI(tie_high_T15Y88), .LO(tie_low_T15Y88));
  sky130_fd_sc_hd__conb_1 conb_T15Y89 (.HI(tie_high_T15Y89), .LO(tie_low_T15Y89));
  sky130_fd_sc_hd__conb_1 conb_T15Y9 (.HI(tie_high_T15Y9), .LO(tie_low_T15Y9));
  sky130_fd_sc_hd__conb_1 conb_T16Y0 (.HI(tie_high_T16Y0), .LO(tie_low_T16Y0));
  sky130_fd_sc_hd__conb_1 conb_T16Y1 (.HI(tie_high_T16Y1), .LO(tie_low_T16Y1));
  sky130_fd_sc_hd__conb_1 conb_T16Y10 (.HI(tie_high_T16Y10), .LO(tie_low_T16Y10));
  sky130_fd_sc_hd__conb_1 conb_T16Y11 (.HI(tie_high_T16Y11), .LO(tie_low_T16Y11));
  sky130_fd_sc_hd__conb_1 conb_T16Y12 (.HI(tie_high_T16Y12), .LO(tie_low_T16Y12));
  sky130_fd_sc_hd__conb_1 conb_T16Y13 (.HI(tie_high_T16Y13), .LO(tie_low_T16Y13));
  sky130_fd_sc_hd__conb_1 conb_T16Y14 (.HI(tie_high_T16Y14), .LO(tie_low_T16Y14));
  sky130_fd_sc_hd__conb_1 conb_T16Y15 (.HI(tie_high_T16Y15), .LO(tie_low_T16Y15));
  sky130_fd_sc_hd__conb_1 conb_T16Y16 (.HI(tie_high_T16Y16), .LO(tie_low_T16Y16));
  sky130_fd_sc_hd__conb_1 conb_T16Y17 (.HI(tie_high_T16Y17), .LO(tie_low_T16Y17));
  sky130_fd_sc_hd__conb_1 conb_T16Y18 (.HI(tie_high_T16Y18), .LO(tie_low_T16Y18));
  sky130_fd_sc_hd__conb_1 conb_T16Y19 (.HI(tie_high_T16Y19), .LO(tie_low_T16Y19));
  sky130_fd_sc_hd__conb_1 conb_T16Y2 (.HI(tie_high_T16Y2), .LO(tie_low_T16Y2));
  sky130_fd_sc_hd__conb_1 conb_T16Y20 (.HI(tie_high_T16Y20), .LO(tie_low_T16Y20));
  sky130_fd_sc_hd__conb_1 conb_T16Y21 (.HI(tie_high_T16Y21), .LO(tie_low_T16Y21));
  sky130_fd_sc_hd__conb_1 conb_T16Y22 (.HI(tie_high_T16Y22), .LO(tie_low_T16Y22));
  sky130_fd_sc_hd__conb_1 conb_T16Y23 (.HI(tie_high_T16Y23), .LO(tie_low_T16Y23));
  sky130_fd_sc_hd__conb_1 conb_T16Y24 (.HI(tie_high_T16Y24), .LO(tie_low_T16Y24));
  sky130_fd_sc_hd__conb_1 conb_T16Y25 (.HI(tie_high_T16Y25), .LO(tie_low_T16Y25));
  sky130_fd_sc_hd__conb_1 conb_T16Y26 (.HI(tie_high_T16Y26), .LO(tie_low_T16Y26));
  sky130_fd_sc_hd__conb_1 conb_T16Y27 (.HI(tie_high_T16Y27), .LO(tie_low_T16Y27));
  sky130_fd_sc_hd__conb_1 conb_T16Y28 (.HI(tie_high_T16Y28), .LO(tie_low_T16Y28));
  sky130_fd_sc_hd__conb_1 conb_T16Y29 (.HI(tie_high_T16Y29), .LO(tie_low_T16Y29));
  sky130_fd_sc_hd__conb_1 conb_T16Y3 (.HI(tie_high_T16Y3), .LO(tie_low_T16Y3));
  sky130_fd_sc_hd__conb_1 conb_T16Y30 (.HI(tie_high_T16Y30), .LO(tie_low_T16Y30));
  sky130_fd_sc_hd__conb_1 conb_T16Y31 (.HI(tie_high_T16Y31), .LO(tie_low_T16Y31));
  sky130_fd_sc_hd__conb_1 conb_T16Y32 (.HI(tie_high_T16Y32), .LO(tie_low_T16Y32));
  sky130_fd_sc_hd__conb_1 conb_T16Y33 (.HI(tie_high_T16Y33), .LO(tie_low_T16Y33));
  sky130_fd_sc_hd__conb_1 conb_T16Y34 (.HI(tie_high_T16Y34), .LO(tie_low_T16Y34));
  sky130_fd_sc_hd__conb_1 conb_T16Y35 (.HI(tie_high_T16Y35), .LO(tie_low_T16Y35));
  sky130_fd_sc_hd__conb_1 conb_T16Y36 (.HI(tie_high_T16Y36), .LO(tie_low_T16Y36));
  sky130_fd_sc_hd__conb_1 conb_T16Y37 (.HI(tie_high_T16Y37), .LO(tie_low_T16Y37));
  sky130_fd_sc_hd__conb_1 conb_T16Y38 (.HI(tie_high_T16Y38), .LO(tie_low_T16Y38));
  sky130_fd_sc_hd__conb_1 conb_T16Y39 (.HI(tie_high_T16Y39), .LO(tie_low_T16Y39));
  sky130_fd_sc_hd__conb_1 conb_T16Y4 (.HI(tie_high_T16Y4), .LO(tie_low_T16Y4));
  sky130_fd_sc_hd__conb_1 conb_T16Y40 (.HI(tie_high_T16Y40), .LO(tie_low_T16Y40));
  sky130_fd_sc_hd__conb_1 conb_T16Y41 (.HI(tie_high_T16Y41), .LO(tie_low_T16Y41));
  sky130_fd_sc_hd__conb_1 conb_T16Y42 (.HI(tie_high_T16Y42), .LO(tie_low_T16Y42));
  sky130_fd_sc_hd__conb_1 conb_T16Y43 (.HI(tie_high_T16Y43), .LO(tie_low_T16Y43));
  sky130_fd_sc_hd__conb_1 conb_T16Y44 (.HI(tie_high_T16Y44), .LO(tie_low_T16Y44));
  sky130_fd_sc_hd__conb_1 conb_T16Y45 (.HI(tie_high_T16Y45), .LO(tie_low_T16Y45));
  sky130_fd_sc_hd__conb_1 conb_T16Y46 (.HI(tie_high_T16Y46), .LO(tie_low_T16Y46));
  sky130_fd_sc_hd__conb_1 conb_T16Y47 (.HI(tie_high_T16Y47), .LO(tie_low_T16Y47));
  sky130_fd_sc_hd__conb_1 conb_T16Y48 (.HI(tie_high_T16Y48), .LO(tie_low_T16Y48));
  sky130_fd_sc_hd__conb_1 conb_T16Y49 (.HI(tie_high_T16Y49), .LO(tie_low_T16Y49));
  sky130_fd_sc_hd__conb_1 conb_T16Y5 (.HI(tie_high_T16Y5), .LO(tie_low_T16Y5));
  sky130_fd_sc_hd__conb_1 conb_T16Y50 (.HI(tie_high_T16Y50), .LO(tie_low_T16Y50));
  sky130_fd_sc_hd__conb_1 conb_T16Y51 (.HI(tie_high_T16Y51), .LO(tie_low_T16Y51));
  sky130_fd_sc_hd__conb_1 conb_T16Y52 (.HI(tie_high_T16Y52), .LO(tie_low_T16Y52));
  sky130_fd_sc_hd__conb_1 conb_T16Y53 (.HI(tie_high_T16Y53), .LO(tie_low_T16Y53));
  sky130_fd_sc_hd__conb_1 conb_T16Y54 (.HI(tie_high_T16Y54), .LO(tie_low_T16Y54));
  sky130_fd_sc_hd__conb_1 conb_T16Y55 (.HI(tie_high_T16Y55), .LO(tie_low_T16Y55));
  sky130_fd_sc_hd__conb_1 conb_T16Y56 (.HI(tie_high_T16Y56), .LO(tie_low_T16Y56));
  sky130_fd_sc_hd__conb_1 conb_T16Y57 (.HI(tie_high_T16Y57), .LO(tie_low_T16Y57));
  sky130_fd_sc_hd__conb_1 conb_T16Y58 (.HI(tie_high_T16Y58), .LO(tie_low_T16Y58));
  sky130_fd_sc_hd__conb_1 conb_T16Y59 (.HI(tie_high_T16Y59), .LO(tie_low_T16Y59));
  sky130_fd_sc_hd__conb_1 conb_T16Y6 (.HI(tie_high_T16Y6), .LO(tie_low_T16Y6));
  sky130_fd_sc_hd__conb_1 conb_T16Y60 (.HI(tie_high_T16Y60), .LO(tie_low_T16Y60));
  sky130_fd_sc_hd__conb_1 conb_T16Y61 (.HI(tie_high_T16Y61), .LO(tie_low_T16Y61));
  sky130_fd_sc_hd__conb_1 conb_T16Y62 (.HI(tie_high_T16Y62), .LO(tie_low_T16Y62));
  sky130_fd_sc_hd__conb_1 conb_T16Y63 (.HI(tie_high_T16Y63), .LO(tie_low_T16Y63));
  sky130_fd_sc_hd__conb_1 conb_T16Y64 (.HI(tie_high_T16Y64), .LO(tie_low_T16Y64));
  sky130_fd_sc_hd__conb_1 conb_T16Y65 (.HI(tie_high_T16Y65), .LO(tie_low_T16Y65));
  sky130_fd_sc_hd__conb_1 conb_T16Y66 (.HI(tie_high_T16Y66), .LO(tie_low_T16Y66));
  sky130_fd_sc_hd__conb_1 conb_T16Y67 (.HI(tie_high_T16Y67), .LO(tie_low_T16Y67));
  sky130_fd_sc_hd__conb_1 conb_T16Y68 (.HI(tie_high_T16Y68), .LO(tie_low_T16Y68));
  sky130_fd_sc_hd__conb_1 conb_T16Y69 (.HI(tie_high_T16Y69), .LO(tie_low_T16Y69));
  sky130_fd_sc_hd__conb_1 conb_T16Y7 (.HI(tie_high_T16Y7), .LO(tie_low_T16Y7));
  sky130_fd_sc_hd__conb_1 conb_T16Y70 (.HI(tie_high_T16Y70), .LO(tie_low_T16Y70));
  sky130_fd_sc_hd__conb_1 conb_T16Y71 (.HI(tie_high_T16Y71), .LO(tie_low_T16Y71));
  sky130_fd_sc_hd__conb_1 conb_T16Y72 (.HI(tie_high_T16Y72), .LO(tie_low_T16Y72));
  sky130_fd_sc_hd__conb_1 conb_T16Y73 (.HI(tie_high_T16Y73), .LO(tie_low_T16Y73));
  sky130_fd_sc_hd__conb_1 conb_T16Y74 (.HI(tie_high_T16Y74), .LO(tie_low_T16Y74));
  sky130_fd_sc_hd__conb_1 conb_T16Y75 (.HI(tie_high_T16Y75), .LO(tie_low_T16Y75));
  sky130_fd_sc_hd__conb_1 conb_T16Y76 (.HI(tie_high_T16Y76), .LO(tie_low_T16Y76));
  sky130_fd_sc_hd__conb_1 conb_T16Y77 (.HI(tie_high_T16Y77), .LO(tie_low_T16Y77));
  sky130_fd_sc_hd__conb_1 conb_T16Y78 (.HI(tie_high_T16Y78), .LO(tie_low_T16Y78));
  sky130_fd_sc_hd__conb_1 conb_T16Y79 (.HI(tie_high_T16Y79), .LO(tie_low_T16Y79));
  sky130_fd_sc_hd__conb_1 conb_T16Y8 (.HI(tie_high_T16Y8), .LO(tie_low_T16Y8));
  sky130_fd_sc_hd__conb_1 conb_T16Y80 (.HI(tie_high_T16Y80), .LO(tie_low_T16Y80));
  sky130_fd_sc_hd__conb_1 conb_T16Y81 (.HI(tie_high_T16Y81), .LO(tie_low_T16Y81));
  sky130_fd_sc_hd__conb_1 conb_T16Y82 (.HI(tie_high_T16Y82), .LO(tie_low_T16Y82));
  sky130_fd_sc_hd__conb_1 conb_T16Y83 (.HI(tie_high_T16Y83), .LO(tie_low_T16Y83));
  sky130_fd_sc_hd__conb_1 conb_T16Y84 (.HI(tie_high_T16Y84), .LO(tie_low_T16Y84));
  sky130_fd_sc_hd__conb_1 conb_T16Y85 (.HI(tie_high_T16Y85), .LO(tie_low_T16Y85));
  sky130_fd_sc_hd__conb_1 conb_T16Y86 (.HI(tie_high_T16Y86), .LO(tie_low_T16Y86));
  sky130_fd_sc_hd__conb_1 conb_T16Y87 (.HI(tie_high_T16Y87), .LO(tie_low_T16Y87));
  sky130_fd_sc_hd__conb_1 conb_T16Y88 (.HI(tie_high_T16Y88), .LO(tie_low_T16Y88));
  sky130_fd_sc_hd__conb_1 conb_T16Y89 (.HI(tie_high_T16Y89), .LO(tie_low_T16Y89));
  sky130_fd_sc_hd__conb_1 conb_T16Y9 (.HI(tie_high_T16Y9), .LO(tie_low_T16Y9));
  sky130_fd_sc_hd__conb_1 conb_T17Y0 (.HI(tie_high_T17Y0), .LO(tie_low_T17Y0));
  sky130_fd_sc_hd__conb_1 conb_T17Y1 (.HI(tie_high_T17Y1), .LO(tie_low_T17Y1));
  sky130_fd_sc_hd__conb_1 conb_T17Y10 (.HI(tie_high_T17Y10), .LO(tie_low_T17Y10));
  sky130_fd_sc_hd__conb_1 conb_T17Y11 (.HI(tie_high_T17Y11), .LO(tie_low_T17Y11));
  sky130_fd_sc_hd__conb_1 conb_T17Y12 (.HI(tie_high_T17Y12), .LO(tie_low_T17Y12));
  sky130_fd_sc_hd__conb_1 conb_T17Y13 (.HI(tie_high_T17Y13), .LO(tie_low_T17Y13));
  sky130_fd_sc_hd__conb_1 conb_T17Y14 (.HI(tie_high_T17Y14), .LO(tie_low_T17Y14));
  sky130_fd_sc_hd__conb_1 conb_T17Y15 (.HI(tie_high_T17Y15), .LO(tie_low_T17Y15));
  sky130_fd_sc_hd__conb_1 conb_T17Y16 (.HI(tie_high_T17Y16), .LO(tie_low_T17Y16));
  sky130_fd_sc_hd__conb_1 conb_T17Y17 (.HI(tie_high_T17Y17), .LO(tie_low_T17Y17));
  sky130_fd_sc_hd__conb_1 conb_T17Y18 (.HI(tie_high_T17Y18), .LO(tie_low_T17Y18));
  sky130_fd_sc_hd__conb_1 conb_T17Y19 (.HI(tie_high_T17Y19), .LO(tie_low_T17Y19));
  sky130_fd_sc_hd__conb_1 conb_T17Y2 (.HI(tie_high_T17Y2), .LO(tie_low_T17Y2));
  sky130_fd_sc_hd__conb_1 conb_T17Y20 (.HI(tie_high_T17Y20), .LO(tie_low_T17Y20));
  sky130_fd_sc_hd__conb_1 conb_T17Y21 (.HI(tie_high_T17Y21), .LO(tie_low_T17Y21));
  sky130_fd_sc_hd__conb_1 conb_T17Y22 (.HI(tie_high_T17Y22), .LO(tie_low_T17Y22));
  sky130_fd_sc_hd__conb_1 conb_T17Y23 (.HI(tie_high_T17Y23), .LO(tie_low_T17Y23));
  sky130_fd_sc_hd__conb_1 conb_T17Y24 (.HI(tie_high_T17Y24), .LO(tie_low_T17Y24));
  sky130_fd_sc_hd__conb_1 conb_T17Y25 (.HI(tie_high_T17Y25), .LO(tie_low_T17Y25));
  sky130_fd_sc_hd__conb_1 conb_T17Y26 (.HI(tie_high_T17Y26), .LO(tie_low_T17Y26));
  sky130_fd_sc_hd__conb_1 conb_T17Y27 (.HI(tie_high_T17Y27), .LO(tie_low_T17Y27));
  sky130_fd_sc_hd__conb_1 conb_T17Y28 (.HI(tie_high_T17Y28), .LO(tie_low_T17Y28));
  sky130_fd_sc_hd__conb_1 conb_T17Y29 (.HI(tie_high_T17Y29), .LO(tie_low_T17Y29));
  sky130_fd_sc_hd__conb_1 conb_T17Y3 (.HI(tie_high_T17Y3), .LO(tie_low_T17Y3));
  sky130_fd_sc_hd__conb_1 conb_T17Y30 (.HI(tie_high_T17Y30), .LO(tie_low_T17Y30));
  sky130_fd_sc_hd__conb_1 conb_T17Y31 (.HI(tie_high_T17Y31), .LO(tie_low_T17Y31));
  sky130_fd_sc_hd__conb_1 conb_T17Y32 (.HI(tie_high_T17Y32), .LO(tie_low_T17Y32));
  sky130_fd_sc_hd__conb_1 conb_T17Y33 (.HI(tie_high_T17Y33), .LO(tie_low_T17Y33));
  sky130_fd_sc_hd__conb_1 conb_T17Y34 (.HI(tie_high_T17Y34), .LO(tie_low_T17Y34));
  sky130_fd_sc_hd__conb_1 conb_T17Y35 (.HI(tie_high_T17Y35), .LO(tie_low_T17Y35));
  sky130_fd_sc_hd__conb_1 conb_T17Y36 (.HI(tie_high_T17Y36), .LO(tie_low_T17Y36));
  sky130_fd_sc_hd__conb_1 conb_T17Y37 (.HI(tie_high_T17Y37), .LO(tie_low_T17Y37));
  sky130_fd_sc_hd__conb_1 conb_T17Y38 (.HI(tie_high_T17Y38), .LO(tie_low_T17Y38));
  sky130_fd_sc_hd__conb_1 conb_T17Y39 (.HI(tie_high_T17Y39), .LO(tie_low_T17Y39));
  sky130_fd_sc_hd__conb_1 conb_T17Y4 (.HI(tie_high_T17Y4), .LO(tie_low_T17Y4));
  sky130_fd_sc_hd__conb_1 conb_T17Y40 (.HI(tie_high_T17Y40), .LO(tie_low_T17Y40));
  sky130_fd_sc_hd__conb_1 conb_T17Y41 (.HI(tie_high_T17Y41), .LO(tie_low_T17Y41));
  sky130_fd_sc_hd__conb_1 conb_T17Y42 (.HI(tie_high_T17Y42), .LO(tie_low_T17Y42));
  sky130_fd_sc_hd__conb_1 conb_T17Y43 (.HI(tie_high_T17Y43), .LO(tie_low_T17Y43));
  sky130_fd_sc_hd__conb_1 conb_T17Y44 (.HI(tie_high_T17Y44), .LO(tie_low_T17Y44));
  sky130_fd_sc_hd__conb_1 conb_T17Y45 (.HI(tie_high_T17Y45), .LO(tie_low_T17Y45));
  sky130_fd_sc_hd__conb_1 conb_T17Y46 (.HI(tie_high_T17Y46), .LO(tie_low_T17Y46));
  sky130_fd_sc_hd__conb_1 conb_T17Y47 (.HI(tie_high_T17Y47), .LO(tie_low_T17Y47));
  sky130_fd_sc_hd__conb_1 conb_T17Y48 (.HI(tie_high_T17Y48), .LO(tie_low_T17Y48));
  sky130_fd_sc_hd__conb_1 conb_T17Y49 (.HI(tie_high_T17Y49), .LO(tie_low_T17Y49));
  sky130_fd_sc_hd__conb_1 conb_T17Y5 (.HI(tie_high_T17Y5), .LO(tie_low_T17Y5));
  sky130_fd_sc_hd__conb_1 conb_T17Y50 (.HI(tie_high_T17Y50), .LO(tie_low_T17Y50));
  sky130_fd_sc_hd__conb_1 conb_T17Y51 (.HI(tie_high_T17Y51), .LO(tie_low_T17Y51));
  sky130_fd_sc_hd__conb_1 conb_T17Y52 (.HI(tie_high_T17Y52), .LO(tie_low_T17Y52));
  sky130_fd_sc_hd__conb_1 conb_T17Y53 (.HI(tie_high_T17Y53), .LO(tie_low_T17Y53));
  sky130_fd_sc_hd__conb_1 conb_T17Y54 (.HI(tie_high_T17Y54), .LO(tie_low_T17Y54));
  sky130_fd_sc_hd__conb_1 conb_T17Y55 (.HI(tie_high_T17Y55), .LO(tie_low_T17Y55));
  sky130_fd_sc_hd__conb_1 conb_T17Y56 (.HI(tie_high_T17Y56), .LO(tie_low_T17Y56));
  sky130_fd_sc_hd__conb_1 conb_T17Y57 (.HI(tie_high_T17Y57), .LO(tie_low_T17Y57));
  sky130_fd_sc_hd__conb_1 conb_T17Y58 (.HI(tie_high_T17Y58), .LO(tie_low_T17Y58));
  sky130_fd_sc_hd__conb_1 conb_T17Y59 (.HI(tie_high_T17Y59), .LO(tie_low_T17Y59));
  sky130_fd_sc_hd__conb_1 conb_T17Y6 (.HI(tie_high_T17Y6), .LO(tie_low_T17Y6));
  sky130_fd_sc_hd__conb_1 conb_T17Y60 (.HI(tie_high_T17Y60), .LO(tie_low_T17Y60));
  sky130_fd_sc_hd__conb_1 conb_T17Y61 (.HI(tie_high_T17Y61), .LO(tie_low_T17Y61));
  sky130_fd_sc_hd__conb_1 conb_T17Y62 (.HI(tie_high_T17Y62), .LO(tie_low_T17Y62));
  sky130_fd_sc_hd__conb_1 conb_T17Y63 (.HI(tie_high_T17Y63), .LO(tie_low_T17Y63));
  sky130_fd_sc_hd__conb_1 conb_T17Y64 (.HI(tie_high_T17Y64), .LO(tie_low_T17Y64));
  sky130_fd_sc_hd__conb_1 conb_T17Y65 (.HI(tie_high_T17Y65), .LO(tie_low_T17Y65));
  sky130_fd_sc_hd__conb_1 conb_T17Y66 (.HI(tie_high_T17Y66), .LO(tie_low_T17Y66));
  sky130_fd_sc_hd__conb_1 conb_T17Y67 (.HI(tie_high_T17Y67), .LO(tie_low_T17Y67));
  sky130_fd_sc_hd__conb_1 conb_T17Y68 (.HI(tie_high_T17Y68), .LO(tie_low_T17Y68));
  sky130_fd_sc_hd__conb_1 conb_T17Y69 (.HI(tie_high_T17Y69), .LO(tie_low_T17Y69));
  sky130_fd_sc_hd__conb_1 conb_T17Y7 (.HI(tie_high_T17Y7), .LO(tie_low_T17Y7));
  sky130_fd_sc_hd__conb_1 conb_T17Y70 (.HI(tie_high_T17Y70), .LO(tie_low_T17Y70));
  sky130_fd_sc_hd__conb_1 conb_T17Y71 (.HI(tie_high_T17Y71), .LO(tie_low_T17Y71));
  sky130_fd_sc_hd__conb_1 conb_T17Y72 (.HI(tie_high_T17Y72), .LO(tie_low_T17Y72));
  sky130_fd_sc_hd__conb_1 conb_T17Y73 (.HI(tie_high_T17Y73), .LO(tie_low_T17Y73));
  sky130_fd_sc_hd__conb_1 conb_T17Y74 (.HI(tie_high_T17Y74), .LO(tie_low_T17Y74));
  sky130_fd_sc_hd__conb_1 conb_T17Y75 (.HI(tie_high_T17Y75), .LO(tie_low_T17Y75));
  sky130_fd_sc_hd__conb_1 conb_T17Y76 (.HI(tie_high_T17Y76), .LO(tie_low_T17Y76));
  sky130_fd_sc_hd__conb_1 conb_T17Y77 (.HI(tie_high_T17Y77), .LO(tie_low_T17Y77));
  sky130_fd_sc_hd__conb_1 conb_T17Y78 (.HI(tie_high_T17Y78), .LO(tie_low_T17Y78));
  sky130_fd_sc_hd__conb_1 conb_T17Y79 (.HI(tie_high_T17Y79), .LO(tie_low_T17Y79));
  sky130_fd_sc_hd__conb_1 conb_T17Y8 (.HI(tie_high_T17Y8), .LO(tie_low_T17Y8));
  sky130_fd_sc_hd__conb_1 conb_T17Y80 (.HI(tie_high_T17Y80), .LO(tie_low_T17Y80));
  sky130_fd_sc_hd__conb_1 conb_T17Y81 (.HI(tie_high_T17Y81), .LO(tie_low_T17Y81));
  sky130_fd_sc_hd__conb_1 conb_T17Y82 (.HI(tie_high_T17Y82), .LO(tie_low_T17Y82));
  sky130_fd_sc_hd__conb_1 conb_T17Y83 (.HI(tie_high_T17Y83), .LO(tie_low_T17Y83));
  sky130_fd_sc_hd__conb_1 conb_T17Y84 (.HI(tie_high_T17Y84), .LO(tie_low_T17Y84));
  sky130_fd_sc_hd__conb_1 conb_T17Y85 (.HI(tie_high_T17Y85), .LO(tie_low_T17Y85));
  sky130_fd_sc_hd__conb_1 conb_T17Y86 (.HI(tie_high_T17Y86), .LO(tie_low_T17Y86));
  sky130_fd_sc_hd__conb_1 conb_T17Y87 (.HI(tie_high_T17Y87), .LO(tie_low_T17Y87));
  sky130_fd_sc_hd__conb_1 conb_T17Y88 (.HI(tie_high_T17Y88), .LO(tie_low_T17Y88));
  sky130_fd_sc_hd__conb_1 conb_T17Y89 (.HI(tie_high_T17Y89), .LO(tie_low_T17Y89));
  sky130_fd_sc_hd__conb_1 conb_T17Y9 (.HI(tie_high_T17Y9), .LO(tie_low_T17Y9));
  sky130_fd_sc_hd__conb_1 conb_T18Y0 (.HI(tie_high_T18Y0), .LO(tie_low_T18Y0));
  sky130_fd_sc_hd__conb_1 conb_T18Y1 (.HI(tie_high_T18Y1), .LO(tie_low_T18Y1));
  sky130_fd_sc_hd__conb_1 conb_T18Y10 (.HI(tie_high_T18Y10), .LO(tie_low_T18Y10));
  sky130_fd_sc_hd__conb_1 conb_T18Y11 (.HI(tie_high_T18Y11), .LO(tie_low_T18Y11));
  sky130_fd_sc_hd__conb_1 conb_T18Y12 (.HI(tie_high_T18Y12), .LO(tie_low_T18Y12));
  sky130_fd_sc_hd__conb_1 conb_T18Y13 (.HI(tie_high_T18Y13), .LO(tie_low_T18Y13));
  sky130_fd_sc_hd__conb_1 conb_T18Y14 (.HI(tie_high_T18Y14), .LO(tie_low_T18Y14));
  sky130_fd_sc_hd__conb_1 conb_T18Y15 (.HI(tie_high_T18Y15), .LO(tie_low_T18Y15));
  sky130_fd_sc_hd__conb_1 conb_T18Y16 (.HI(tie_high_T18Y16), .LO(tie_low_T18Y16));
  sky130_fd_sc_hd__conb_1 conb_T18Y17 (.HI(tie_high_T18Y17), .LO(tie_low_T18Y17));
  sky130_fd_sc_hd__conb_1 conb_T18Y18 (.HI(tie_high_T18Y18), .LO(tie_low_T18Y18));
  sky130_fd_sc_hd__conb_1 conb_T18Y19 (.HI(tie_high_T18Y19), .LO(tie_low_T18Y19));
  sky130_fd_sc_hd__conb_1 conb_T18Y2 (.HI(tie_high_T18Y2), .LO(tie_low_T18Y2));
  sky130_fd_sc_hd__conb_1 conb_T18Y20 (.HI(tie_high_T18Y20), .LO(tie_low_T18Y20));
  sky130_fd_sc_hd__conb_1 conb_T18Y21 (.HI(tie_high_T18Y21), .LO(tie_low_T18Y21));
  sky130_fd_sc_hd__conb_1 conb_T18Y22 (.HI(tie_high_T18Y22), .LO(tie_low_T18Y22));
  sky130_fd_sc_hd__conb_1 conb_T18Y23 (.HI(tie_high_T18Y23), .LO(tie_low_T18Y23));
  sky130_fd_sc_hd__conb_1 conb_T18Y24 (.HI(tie_high_T18Y24), .LO(tie_low_T18Y24));
  sky130_fd_sc_hd__conb_1 conb_T18Y25 (.HI(tie_high_T18Y25), .LO(tie_low_T18Y25));
  sky130_fd_sc_hd__conb_1 conb_T18Y26 (.HI(tie_high_T18Y26), .LO(tie_low_T18Y26));
  sky130_fd_sc_hd__conb_1 conb_T18Y27 (.HI(tie_high_T18Y27), .LO(tie_low_T18Y27));
  sky130_fd_sc_hd__conb_1 conb_T18Y28 (.HI(tie_high_T18Y28), .LO(tie_low_T18Y28));
  sky130_fd_sc_hd__conb_1 conb_T18Y29 (.HI(tie_high_T18Y29), .LO(tie_low_T18Y29));
  sky130_fd_sc_hd__conb_1 conb_T18Y3 (.HI(tie_high_T18Y3), .LO(tie_low_T18Y3));
  sky130_fd_sc_hd__conb_1 conb_T18Y30 (.HI(tie_high_T18Y30), .LO(tie_low_T18Y30));
  sky130_fd_sc_hd__conb_1 conb_T18Y31 (.HI(tie_high_T18Y31), .LO(tie_low_T18Y31));
  sky130_fd_sc_hd__conb_1 conb_T18Y32 (.HI(tie_high_T18Y32), .LO(tie_low_T18Y32));
  sky130_fd_sc_hd__conb_1 conb_T18Y33 (.HI(tie_high_T18Y33), .LO(tie_low_T18Y33));
  sky130_fd_sc_hd__conb_1 conb_T18Y34 (.HI(tie_high_T18Y34), .LO(tie_low_T18Y34));
  sky130_fd_sc_hd__conb_1 conb_T18Y35 (.HI(tie_high_T18Y35), .LO(tie_low_T18Y35));
  sky130_fd_sc_hd__conb_1 conb_T18Y36 (.HI(tie_high_T18Y36), .LO(tie_low_T18Y36));
  sky130_fd_sc_hd__conb_1 conb_T18Y37 (.HI(tie_high_T18Y37), .LO(tie_low_T18Y37));
  sky130_fd_sc_hd__conb_1 conb_T18Y38 (.HI(tie_high_T18Y38), .LO(tie_low_T18Y38));
  sky130_fd_sc_hd__conb_1 conb_T18Y39 (.HI(tie_high_T18Y39), .LO(tie_low_T18Y39));
  sky130_fd_sc_hd__conb_1 conb_T18Y4 (.HI(tie_high_T18Y4), .LO(tie_low_T18Y4));
  sky130_fd_sc_hd__conb_1 conb_T18Y40 (.HI(tie_high_T18Y40), .LO(tie_low_T18Y40));
  sky130_fd_sc_hd__conb_1 conb_T18Y41 (.HI(tie_high_T18Y41), .LO(tie_low_T18Y41));
  sky130_fd_sc_hd__conb_1 conb_T18Y42 (.HI(tie_high_T18Y42), .LO(tie_low_T18Y42));
  sky130_fd_sc_hd__conb_1 conb_T18Y43 (.HI(tie_high_T18Y43), .LO(tie_low_T18Y43));
  sky130_fd_sc_hd__conb_1 conb_T18Y44 (.HI(tie_high_T18Y44), .LO(tie_low_T18Y44));
  sky130_fd_sc_hd__conb_1 conb_T18Y45 (.HI(tie_high_T18Y45), .LO(tie_low_T18Y45));
  sky130_fd_sc_hd__conb_1 conb_T18Y46 (.HI(tie_high_T18Y46), .LO(tie_low_T18Y46));
  sky130_fd_sc_hd__conb_1 conb_T18Y47 (.HI(tie_high_T18Y47), .LO(tie_low_T18Y47));
  sky130_fd_sc_hd__conb_1 conb_T18Y48 (.HI(tie_high_T18Y48), .LO(tie_low_T18Y48));
  sky130_fd_sc_hd__conb_1 conb_T18Y49 (.HI(tie_high_T18Y49), .LO(tie_low_T18Y49));
  sky130_fd_sc_hd__conb_1 conb_T18Y5 (.HI(tie_high_T18Y5), .LO(tie_low_T18Y5));
  sky130_fd_sc_hd__conb_1 conb_T18Y50 (.HI(tie_high_T18Y50), .LO(tie_low_T18Y50));
  sky130_fd_sc_hd__conb_1 conb_T18Y51 (.HI(tie_high_T18Y51), .LO(tie_low_T18Y51));
  sky130_fd_sc_hd__conb_1 conb_T18Y52 (.HI(tie_high_T18Y52), .LO(tie_low_T18Y52));
  sky130_fd_sc_hd__conb_1 conb_T18Y53 (.HI(tie_high_T18Y53), .LO(tie_low_T18Y53));
  sky130_fd_sc_hd__conb_1 conb_T18Y54 (.HI(tie_high_T18Y54), .LO(tie_low_T18Y54));
  sky130_fd_sc_hd__conb_1 conb_T18Y55 (.HI(tie_high_T18Y55), .LO(tie_low_T18Y55));
  sky130_fd_sc_hd__conb_1 conb_T18Y56 (.HI(tie_high_T18Y56), .LO(tie_low_T18Y56));
  sky130_fd_sc_hd__conb_1 conb_T18Y57 (.HI(tie_high_T18Y57), .LO(tie_low_T18Y57));
  sky130_fd_sc_hd__conb_1 conb_T18Y58 (.HI(tie_high_T18Y58), .LO(tie_low_T18Y58));
  sky130_fd_sc_hd__conb_1 conb_T18Y59 (.HI(tie_high_T18Y59), .LO(tie_low_T18Y59));
  sky130_fd_sc_hd__conb_1 conb_T18Y6 (.HI(tie_high_T18Y6), .LO(tie_low_T18Y6));
  sky130_fd_sc_hd__conb_1 conb_T18Y60 (.HI(tie_high_T18Y60), .LO(tie_low_T18Y60));
  sky130_fd_sc_hd__conb_1 conb_T18Y61 (.HI(tie_high_T18Y61), .LO(tie_low_T18Y61));
  sky130_fd_sc_hd__conb_1 conb_T18Y62 (.HI(tie_high_T18Y62), .LO(tie_low_T18Y62));
  sky130_fd_sc_hd__conb_1 conb_T18Y63 (.HI(tie_high_T18Y63), .LO(tie_low_T18Y63));
  sky130_fd_sc_hd__conb_1 conb_T18Y64 (.HI(tie_high_T18Y64), .LO(tie_low_T18Y64));
  sky130_fd_sc_hd__conb_1 conb_T18Y65 (.HI(tie_high_T18Y65), .LO(tie_low_T18Y65));
  sky130_fd_sc_hd__conb_1 conb_T18Y66 (.HI(tie_high_T18Y66), .LO(tie_low_T18Y66));
  sky130_fd_sc_hd__conb_1 conb_T18Y67 (.HI(tie_high_T18Y67), .LO(tie_low_T18Y67));
  sky130_fd_sc_hd__conb_1 conb_T18Y68 (.HI(tie_high_T18Y68), .LO(tie_low_T18Y68));
  sky130_fd_sc_hd__conb_1 conb_T18Y69 (.HI(tie_high_T18Y69), .LO(tie_low_T18Y69));
  sky130_fd_sc_hd__conb_1 conb_T18Y7 (.HI(tie_high_T18Y7), .LO(tie_low_T18Y7));
  sky130_fd_sc_hd__conb_1 conb_T18Y70 (.HI(tie_high_T18Y70), .LO(tie_low_T18Y70));
  sky130_fd_sc_hd__conb_1 conb_T18Y71 (.HI(tie_high_T18Y71), .LO(tie_low_T18Y71));
  sky130_fd_sc_hd__conb_1 conb_T18Y72 (.HI(tie_high_T18Y72), .LO(tie_low_T18Y72));
  sky130_fd_sc_hd__conb_1 conb_T18Y73 (.HI(tie_high_T18Y73), .LO(tie_low_T18Y73));
  sky130_fd_sc_hd__conb_1 conb_T18Y74 (.HI(tie_high_T18Y74), .LO(tie_low_T18Y74));
  sky130_fd_sc_hd__conb_1 conb_T18Y75 (.HI(tie_high_T18Y75), .LO(tie_low_T18Y75));
  sky130_fd_sc_hd__conb_1 conb_T18Y76 (.HI(tie_high_T18Y76), .LO(tie_low_T18Y76));
  sky130_fd_sc_hd__conb_1 conb_T18Y77 (.HI(tie_high_T18Y77), .LO(tie_low_T18Y77));
  sky130_fd_sc_hd__conb_1 conb_T18Y78 (.HI(tie_high_T18Y78), .LO(tie_low_T18Y78));
  sky130_fd_sc_hd__conb_1 conb_T18Y79 (.HI(tie_high_T18Y79), .LO(tie_low_T18Y79));
  sky130_fd_sc_hd__conb_1 conb_T18Y8 (.HI(tie_high_T18Y8), .LO(tie_low_T18Y8));
  sky130_fd_sc_hd__conb_1 conb_T18Y80 (.HI(tie_high_T18Y80), .LO(tie_low_T18Y80));
  sky130_fd_sc_hd__conb_1 conb_T18Y81 (.HI(tie_high_T18Y81), .LO(tie_low_T18Y81));
  sky130_fd_sc_hd__conb_1 conb_T18Y82 (.HI(tie_high_T18Y82), .LO(tie_low_T18Y82));
  sky130_fd_sc_hd__conb_1 conb_T18Y83 (.HI(tie_high_T18Y83), .LO(tie_low_T18Y83));
  sky130_fd_sc_hd__conb_1 conb_T18Y84 (.HI(tie_high_T18Y84), .LO(tie_low_T18Y84));
  sky130_fd_sc_hd__conb_1 conb_T18Y85 (.HI(tie_high_T18Y85), .LO(tie_low_T18Y85));
  sky130_fd_sc_hd__conb_1 conb_T18Y86 (.HI(tie_high_T18Y86), .LO(tie_low_T18Y86));
  sky130_fd_sc_hd__conb_1 conb_T18Y87 (.HI(tie_high_T18Y87), .LO(tie_low_T18Y87));
  sky130_fd_sc_hd__conb_1 conb_T18Y88 (.HI(tie_high_T18Y88), .LO(tie_low_T18Y88));
  sky130_fd_sc_hd__conb_1 conb_T18Y89 (.HI(tie_high_T18Y89), .LO(tie_low_T18Y89));
  sky130_fd_sc_hd__conb_1 conb_T18Y9 (.HI(tie_high_T18Y9), .LO(tie_low_T18Y9));
  sky130_fd_sc_hd__conb_1 conb_T19Y0 (.HI(tie_high_T19Y0), .LO(tie_low_T19Y0));
  sky130_fd_sc_hd__conb_1 conb_T19Y1 (.HI(tie_high_T19Y1), .LO(tie_low_T19Y1));
  sky130_fd_sc_hd__conb_1 conb_T19Y10 (.HI(tie_high_T19Y10), .LO(tie_low_T19Y10));
  sky130_fd_sc_hd__conb_1 conb_T19Y11 (.HI(tie_high_T19Y11), .LO(tie_low_T19Y11));
  sky130_fd_sc_hd__conb_1 conb_T19Y12 (.HI(tie_high_T19Y12), .LO(tie_low_T19Y12));
  sky130_fd_sc_hd__conb_1 conb_T19Y13 (.HI(tie_high_T19Y13), .LO(tie_low_T19Y13));
  sky130_fd_sc_hd__conb_1 conb_T19Y14 (.HI(tie_high_T19Y14), .LO(tie_low_T19Y14));
  sky130_fd_sc_hd__conb_1 conb_T19Y15 (.HI(tie_high_T19Y15), .LO(tie_low_T19Y15));
  sky130_fd_sc_hd__conb_1 conb_T19Y16 (.HI(tie_high_T19Y16), .LO(tie_low_T19Y16));
  sky130_fd_sc_hd__conb_1 conb_T19Y17 (.HI(tie_high_T19Y17), .LO(tie_low_T19Y17));
  sky130_fd_sc_hd__conb_1 conb_T19Y18 (.HI(tie_high_T19Y18), .LO(tie_low_T19Y18));
  sky130_fd_sc_hd__conb_1 conb_T19Y19 (.HI(tie_high_T19Y19), .LO(tie_low_T19Y19));
  sky130_fd_sc_hd__conb_1 conb_T19Y2 (.HI(tie_high_T19Y2), .LO(tie_low_T19Y2));
  sky130_fd_sc_hd__conb_1 conb_T19Y20 (.HI(tie_high_T19Y20), .LO(tie_low_T19Y20));
  sky130_fd_sc_hd__conb_1 conb_T19Y21 (.HI(tie_high_T19Y21), .LO(tie_low_T19Y21));
  sky130_fd_sc_hd__conb_1 conb_T19Y22 (.HI(tie_high_T19Y22), .LO(tie_low_T19Y22));
  sky130_fd_sc_hd__conb_1 conb_T19Y23 (.HI(tie_high_T19Y23), .LO(tie_low_T19Y23));
  sky130_fd_sc_hd__conb_1 conb_T19Y24 (.HI(tie_high_T19Y24), .LO(tie_low_T19Y24));
  sky130_fd_sc_hd__conb_1 conb_T19Y25 (.HI(tie_high_T19Y25), .LO(tie_low_T19Y25));
  sky130_fd_sc_hd__conb_1 conb_T19Y26 (.HI(tie_high_T19Y26), .LO(tie_low_T19Y26));
  sky130_fd_sc_hd__conb_1 conb_T19Y27 (.HI(tie_high_T19Y27), .LO(tie_low_T19Y27));
  sky130_fd_sc_hd__conb_1 conb_T19Y28 (.HI(tie_high_T19Y28), .LO(tie_low_T19Y28));
  sky130_fd_sc_hd__conb_1 conb_T19Y29 (.HI(tie_high_T19Y29), .LO(tie_low_T19Y29));
  sky130_fd_sc_hd__conb_1 conb_T19Y3 (.HI(tie_high_T19Y3), .LO(tie_low_T19Y3));
  sky130_fd_sc_hd__conb_1 conb_T19Y30 (.HI(tie_high_T19Y30), .LO(tie_low_T19Y30));
  sky130_fd_sc_hd__conb_1 conb_T19Y31 (.HI(tie_high_T19Y31), .LO(tie_low_T19Y31));
  sky130_fd_sc_hd__conb_1 conb_T19Y32 (.HI(tie_high_T19Y32), .LO(tie_low_T19Y32));
  sky130_fd_sc_hd__conb_1 conb_T19Y33 (.HI(tie_high_T19Y33), .LO(tie_low_T19Y33));
  sky130_fd_sc_hd__conb_1 conb_T19Y34 (.HI(tie_high_T19Y34), .LO(tie_low_T19Y34));
  sky130_fd_sc_hd__conb_1 conb_T19Y35 (.HI(tie_high_T19Y35), .LO(tie_low_T19Y35));
  sky130_fd_sc_hd__conb_1 conb_T19Y36 (.HI(tie_high_T19Y36), .LO(tie_low_T19Y36));
  sky130_fd_sc_hd__conb_1 conb_T19Y37 (.HI(tie_high_T19Y37), .LO(tie_low_T19Y37));
  sky130_fd_sc_hd__conb_1 conb_T19Y38 (.HI(tie_high_T19Y38), .LO(tie_low_T19Y38));
  sky130_fd_sc_hd__conb_1 conb_T19Y39 (.HI(tie_high_T19Y39), .LO(tie_low_T19Y39));
  sky130_fd_sc_hd__conb_1 conb_T19Y4 (.HI(tie_high_T19Y4), .LO(tie_low_T19Y4));
  sky130_fd_sc_hd__conb_1 conb_T19Y40 (.HI(tie_high_T19Y40), .LO(tie_low_T19Y40));
  sky130_fd_sc_hd__conb_1 conb_T19Y41 (.HI(tie_high_T19Y41), .LO(tie_low_T19Y41));
  sky130_fd_sc_hd__conb_1 conb_T19Y42 (.HI(tie_high_T19Y42), .LO(tie_low_T19Y42));
  sky130_fd_sc_hd__conb_1 conb_T19Y43 (.HI(tie_high_T19Y43), .LO(tie_low_T19Y43));
  sky130_fd_sc_hd__conb_1 conb_T19Y44 (.HI(tie_high_T19Y44), .LO(tie_low_T19Y44));
  sky130_fd_sc_hd__conb_1 conb_T19Y45 (.HI(tie_high_T19Y45), .LO(tie_low_T19Y45));
  sky130_fd_sc_hd__conb_1 conb_T19Y46 (.HI(tie_high_T19Y46), .LO(tie_low_T19Y46));
  sky130_fd_sc_hd__conb_1 conb_T19Y47 (.HI(tie_high_T19Y47), .LO(tie_low_T19Y47));
  sky130_fd_sc_hd__conb_1 conb_T19Y48 (.HI(tie_high_T19Y48), .LO(tie_low_T19Y48));
  sky130_fd_sc_hd__conb_1 conb_T19Y49 (.HI(tie_high_T19Y49), .LO(tie_low_T19Y49));
  sky130_fd_sc_hd__conb_1 conb_T19Y5 (.HI(tie_high_T19Y5), .LO(tie_low_T19Y5));
  sky130_fd_sc_hd__conb_1 conb_T19Y50 (.HI(tie_high_T19Y50), .LO(tie_low_T19Y50));
  sky130_fd_sc_hd__conb_1 conb_T19Y51 (.HI(tie_high_T19Y51), .LO(tie_low_T19Y51));
  sky130_fd_sc_hd__conb_1 conb_T19Y52 (.HI(tie_high_T19Y52), .LO(tie_low_T19Y52));
  sky130_fd_sc_hd__conb_1 conb_T19Y53 (.HI(tie_high_T19Y53), .LO(tie_low_T19Y53));
  sky130_fd_sc_hd__conb_1 conb_T19Y54 (.HI(tie_high_T19Y54), .LO(tie_low_T19Y54));
  sky130_fd_sc_hd__conb_1 conb_T19Y55 (.HI(tie_high_T19Y55), .LO(tie_low_T19Y55));
  sky130_fd_sc_hd__conb_1 conb_T19Y56 (.HI(tie_high_T19Y56), .LO(tie_low_T19Y56));
  sky130_fd_sc_hd__conb_1 conb_T19Y57 (.HI(tie_high_T19Y57), .LO(tie_low_T19Y57));
  sky130_fd_sc_hd__conb_1 conb_T19Y58 (.HI(tie_high_T19Y58), .LO(tie_low_T19Y58));
  sky130_fd_sc_hd__conb_1 conb_T19Y59 (.HI(tie_high_T19Y59), .LO(tie_low_T19Y59));
  sky130_fd_sc_hd__conb_1 conb_T19Y6 (.HI(tie_high_T19Y6), .LO(tie_low_T19Y6));
  sky130_fd_sc_hd__conb_1 conb_T19Y60 (.HI(tie_high_T19Y60), .LO(tie_low_T19Y60));
  sky130_fd_sc_hd__conb_1 conb_T19Y61 (.HI(tie_high_T19Y61), .LO(tie_low_T19Y61));
  sky130_fd_sc_hd__conb_1 conb_T19Y62 (.HI(tie_high_T19Y62), .LO(tie_low_T19Y62));
  sky130_fd_sc_hd__conb_1 conb_T19Y63 (.HI(tie_high_T19Y63), .LO(tie_low_T19Y63));
  sky130_fd_sc_hd__conb_1 conb_T19Y64 (.HI(tie_high_T19Y64), .LO(tie_low_T19Y64));
  sky130_fd_sc_hd__conb_1 conb_T19Y65 (.HI(tie_high_T19Y65), .LO(tie_low_T19Y65));
  sky130_fd_sc_hd__conb_1 conb_T19Y66 (.HI(tie_high_T19Y66), .LO(tie_low_T19Y66));
  sky130_fd_sc_hd__conb_1 conb_T19Y67 (.HI(tie_high_T19Y67), .LO(tie_low_T19Y67));
  sky130_fd_sc_hd__conb_1 conb_T19Y68 (.HI(tie_high_T19Y68), .LO(tie_low_T19Y68));
  sky130_fd_sc_hd__conb_1 conb_T19Y69 (.HI(tie_high_T19Y69), .LO(tie_low_T19Y69));
  sky130_fd_sc_hd__conb_1 conb_T19Y7 (.HI(tie_high_T19Y7), .LO(tie_low_T19Y7));
  sky130_fd_sc_hd__conb_1 conb_T19Y70 (.HI(tie_high_T19Y70), .LO(tie_low_T19Y70));
  sky130_fd_sc_hd__conb_1 conb_T19Y71 (.HI(tie_high_T19Y71), .LO(tie_low_T19Y71));
  sky130_fd_sc_hd__conb_1 conb_T19Y72 (.HI(tie_high_T19Y72), .LO(tie_low_T19Y72));
  sky130_fd_sc_hd__conb_1 conb_T19Y73 (.HI(tie_high_T19Y73), .LO(tie_low_T19Y73));
  sky130_fd_sc_hd__conb_1 conb_T19Y74 (.HI(tie_high_T19Y74), .LO(tie_low_T19Y74));
  sky130_fd_sc_hd__conb_1 conb_T19Y75 (.HI(tie_high_T19Y75), .LO(tie_low_T19Y75));
  sky130_fd_sc_hd__conb_1 conb_T19Y76 (.HI(tie_high_T19Y76), .LO(tie_low_T19Y76));
  sky130_fd_sc_hd__conb_1 conb_T19Y77 (.HI(tie_high_T19Y77), .LO(tie_low_T19Y77));
  sky130_fd_sc_hd__conb_1 conb_T19Y78 (.HI(tie_high_T19Y78), .LO(tie_low_T19Y78));
  sky130_fd_sc_hd__conb_1 conb_T19Y79 (.HI(tie_high_T19Y79), .LO(tie_low_T19Y79));
  sky130_fd_sc_hd__conb_1 conb_T19Y8 (.HI(tie_high_T19Y8), .LO(tie_low_T19Y8));
  sky130_fd_sc_hd__conb_1 conb_T19Y80 (.HI(tie_high_T19Y80), .LO(tie_low_T19Y80));
  sky130_fd_sc_hd__conb_1 conb_T19Y81 (.HI(tie_high_T19Y81), .LO(tie_low_T19Y81));
  sky130_fd_sc_hd__conb_1 conb_T19Y82 (.HI(tie_high_T19Y82), .LO(tie_low_T19Y82));
  sky130_fd_sc_hd__conb_1 conb_T19Y83 (.HI(tie_high_T19Y83), .LO(tie_low_T19Y83));
  sky130_fd_sc_hd__conb_1 conb_T19Y84 (.HI(tie_high_T19Y84), .LO(tie_low_T19Y84));
  sky130_fd_sc_hd__conb_1 conb_T19Y85 (.HI(tie_high_T19Y85), .LO(tie_low_T19Y85));
  sky130_fd_sc_hd__conb_1 conb_T19Y86 (.HI(tie_high_T19Y86), .LO(tie_low_T19Y86));
  sky130_fd_sc_hd__conb_1 conb_T19Y87 (.HI(tie_high_T19Y87), .LO(tie_low_T19Y87));
  sky130_fd_sc_hd__conb_1 conb_T19Y88 (.HI(tie_high_T19Y88), .LO(tie_low_T19Y88));
  sky130_fd_sc_hd__conb_1 conb_T19Y89 (.HI(tie_high_T19Y89), .LO(tie_low_T19Y89));
  sky130_fd_sc_hd__conb_1 conb_T19Y9 (.HI(tie_high_T19Y9), .LO(tie_low_T19Y9));
  sky130_fd_sc_hd__conb_1 conb_T1Y0 (.HI(tie_high_T1Y0), .LO(tie_low_T1Y0));
  sky130_fd_sc_hd__conb_1 conb_T1Y1 (.HI(tie_high_T1Y1), .LO(tie_low_T1Y1));
  sky130_fd_sc_hd__conb_1 conb_T1Y10 (.HI(tie_high_T1Y10), .LO(tie_low_T1Y10));
  sky130_fd_sc_hd__conb_1 conb_T1Y11 (.HI(tie_high_T1Y11), .LO(tie_low_T1Y11));
  sky130_fd_sc_hd__conb_1 conb_T1Y12 (.HI(tie_high_T1Y12), .LO(tie_low_T1Y12));
  sky130_fd_sc_hd__conb_1 conb_T1Y13 (.HI(tie_high_T1Y13), .LO(tie_low_T1Y13));
  sky130_fd_sc_hd__conb_1 conb_T1Y14 (.HI(tie_high_T1Y14), .LO(tie_low_T1Y14));
  sky130_fd_sc_hd__conb_1 conb_T1Y15 (.HI(tie_high_T1Y15), .LO(tie_low_T1Y15));
  sky130_fd_sc_hd__conb_1 conb_T1Y16 (.HI(tie_high_T1Y16), .LO(tie_low_T1Y16));
  sky130_fd_sc_hd__conb_1 conb_T1Y17 (.HI(tie_high_T1Y17), .LO(tie_low_T1Y17));
  sky130_fd_sc_hd__conb_1 conb_T1Y18 (.HI(tie_high_T1Y18), .LO(tie_low_T1Y18));
  sky130_fd_sc_hd__conb_1 conb_T1Y19 (.HI(tie_high_T1Y19), .LO(tie_low_T1Y19));
  sky130_fd_sc_hd__conb_1 conb_T1Y2 (.HI(tie_high_T1Y2), .LO(tie_low_T1Y2));
  sky130_fd_sc_hd__conb_1 conb_T1Y20 (.HI(tie_high_T1Y20), .LO(tie_low_T1Y20));
  sky130_fd_sc_hd__conb_1 conb_T1Y21 (.HI(tie_high_T1Y21), .LO(tie_low_T1Y21));
  sky130_fd_sc_hd__conb_1 conb_T1Y22 (.HI(tie_high_T1Y22), .LO(tie_low_T1Y22));
  sky130_fd_sc_hd__conb_1 conb_T1Y23 (.HI(tie_high_T1Y23), .LO(tie_low_T1Y23));
  sky130_fd_sc_hd__conb_1 conb_T1Y24 (.HI(tie_high_T1Y24), .LO(tie_low_T1Y24));
  sky130_fd_sc_hd__conb_1 conb_T1Y25 (.HI(tie_high_T1Y25), .LO(tie_low_T1Y25));
  sky130_fd_sc_hd__conb_1 conb_T1Y26 (.HI(tie_high_T1Y26), .LO(tie_low_T1Y26));
  sky130_fd_sc_hd__conb_1 conb_T1Y27 (.HI(tie_high_T1Y27), .LO(tie_low_T1Y27));
  sky130_fd_sc_hd__conb_1 conb_T1Y28 (.HI(tie_high_T1Y28), .LO(tie_low_T1Y28));
  sky130_fd_sc_hd__conb_1 conb_T1Y29 (.HI(tie_high_T1Y29), .LO(tie_low_T1Y29));
  sky130_fd_sc_hd__conb_1 conb_T1Y3 (.HI(tie_high_T1Y3), .LO(tie_low_T1Y3));
  sky130_fd_sc_hd__conb_1 conb_T1Y30 (.HI(tie_high_T1Y30), .LO(tie_low_T1Y30));
  sky130_fd_sc_hd__conb_1 conb_T1Y31 (.HI(tie_high_T1Y31), .LO(tie_low_T1Y31));
  sky130_fd_sc_hd__conb_1 conb_T1Y32 (.HI(tie_high_T1Y32), .LO(tie_low_T1Y32));
  sky130_fd_sc_hd__conb_1 conb_T1Y33 (.HI(tie_high_T1Y33), .LO(tie_low_T1Y33));
  sky130_fd_sc_hd__conb_1 conb_T1Y34 (.HI(tie_high_T1Y34), .LO(tie_low_T1Y34));
  sky130_fd_sc_hd__conb_1 conb_T1Y35 (.HI(tie_high_T1Y35), .LO(tie_low_T1Y35));
  sky130_fd_sc_hd__conb_1 conb_T1Y36 (.HI(tie_high_T1Y36), .LO(tie_low_T1Y36));
  sky130_fd_sc_hd__conb_1 conb_T1Y37 (.HI(tie_high_T1Y37), .LO(tie_low_T1Y37));
  sky130_fd_sc_hd__conb_1 conb_T1Y38 (.HI(tie_high_T1Y38), .LO(tie_low_T1Y38));
  sky130_fd_sc_hd__conb_1 conb_T1Y39 (.HI(tie_high_T1Y39), .LO(tie_low_T1Y39));
  sky130_fd_sc_hd__conb_1 conb_T1Y4 (.HI(tie_high_T1Y4), .LO(tie_low_T1Y4));
  sky130_fd_sc_hd__conb_1 conb_T1Y40 (.HI(tie_high_T1Y40), .LO(tie_low_T1Y40));
  sky130_fd_sc_hd__conb_1 conb_T1Y41 (.HI(tie_high_T1Y41), .LO(tie_low_T1Y41));
  sky130_fd_sc_hd__conb_1 conb_T1Y42 (.HI(tie_high_T1Y42), .LO(tie_low_T1Y42));
  sky130_fd_sc_hd__conb_1 conb_T1Y43 (.HI(tie_high_T1Y43), .LO(tie_low_T1Y43));
  sky130_fd_sc_hd__conb_1 conb_T1Y44 (.HI(tie_high_T1Y44), .LO(tie_low_T1Y44));
  sky130_fd_sc_hd__conb_1 conb_T1Y45 (.HI(tie_high_T1Y45), .LO(tie_low_T1Y45));
  sky130_fd_sc_hd__conb_1 conb_T1Y46 (.HI(tie_high_T1Y46), .LO(tie_low_T1Y46));
  sky130_fd_sc_hd__conb_1 conb_T1Y47 (.HI(tie_high_T1Y47), .LO(tie_low_T1Y47));
  sky130_fd_sc_hd__conb_1 conb_T1Y48 (.HI(tie_high_T1Y48), .LO(tie_low_T1Y48));
  sky130_fd_sc_hd__conb_1 conb_T1Y49 (.HI(tie_high_T1Y49), .LO(tie_low_T1Y49));
  sky130_fd_sc_hd__conb_1 conb_T1Y5 (.HI(tie_high_T1Y5), .LO(tie_low_T1Y5));
  sky130_fd_sc_hd__conb_1 conb_T1Y50 (.HI(tie_high_T1Y50), .LO(tie_low_T1Y50));
  sky130_fd_sc_hd__conb_1 conb_T1Y51 (.HI(tie_high_T1Y51), .LO(tie_low_T1Y51));
  sky130_fd_sc_hd__conb_1 conb_T1Y52 (.HI(tie_high_T1Y52), .LO(tie_low_T1Y52));
  sky130_fd_sc_hd__conb_1 conb_T1Y53 (.HI(tie_high_T1Y53), .LO(tie_low_T1Y53));
  sky130_fd_sc_hd__conb_1 conb_T1Y54 (.HI(tie_high_T1Y54), .LO(tie_low_T1Y54));
  sky130_fd_sc_hd__conb_1 conb_T1Y55 (.HI(tie_high_T1Y55), .LO(tie_low_T1Y55));
  sky130_fd_sc_hd__conb_1 conb_T1Y56 (.HI(tie_high_T1Y56), .LO(tie_low_T1Y56));
  sky130_fd_sc_hd__conb_1 conb_T1Y57 (.HI(tie_high_T1Y57), .LO(tie_low_T1Y57));
  sky130_fd_sc_hd__conb_1 conb_T1Y58 (.HI(tie_high_T1Y58), .LO(tie_low_T1Y58));
  sky130_fd_sc_hd__conb_1 conb_T1Y59 (.HI(tie_high_T1Y59), .LO(tie_low_T1Y59));
  sky130_fd_sc_hd__conb_1 conb_T1Y6 (.HI(tie_high_T1Y6), .LO(tie_low_T1Y6));
  sky130_fd_sc_hd__conb_1 conb_T1Y60 (.HI(tie_high_T1Y60), .LO(tie_low_T1Y60));
  sky130_fd_sc_hd__conb_1 conb_T1Y61 (.HI(tie_high_T1Y61), .LO(tie_low_T1Y61));
  sky130_fd_sc_hd__conb_1 conb_T1Y62 (.HI(tie_high_T1Y62), .LO(tie_low_T1Y62));
  sky130_fd_sc_hd__conb_1 conb_T1Y63 (.HI(tie_high_T1Y63), .LO(tie_low_T1Y63));
  sky130_fd_sc_hd__conb_1 conb_T1Y64 (.HI(tie_high_T1Y64), .LO(tie_low_T1Y64));
  sky130_fd_sc_hd__conb_1 conb_T1Y65 (.HI(tie_high_T1Y65), .LO(tie_low_T1Y65));
  sky130_fd_sc_hd__conb_1 conb_T1Y66 (.HI(tie_high_T1Y66), .LO(tie_low_T1Y66));
  sky130_fd_sc_hd__conb_1 conb_T1Y67 (.HI(tie_high_T1Y67), .LO(tie_low_T1Y67));
  sky130_fd_sc_hd__conb_1 conb_T1Y68 (.HI(tie_high_T1Y68), .LO(tie_low_T1Y68));
  sky130_fd_sc_hd__conb_1 conb_T1Y69 (.HI(tie_high_T1Y69), .LO(tie_low_T1Y69));
  sky130_fd_sc_hd__conb_1 conb_T1Y7 (.HI(tie_high_T1Y7), .LO(tie_low_T1Y7));
  sky130_fd_sc_hd__conb_1 conb_T1Y70 (.HI(tie_high_T1Y70), .LO(tie_low_T1Y70));
  sky130_fd_sc_hd__conb_1 conb_T1Y71 (.HI(tie_high_T1Y71), .LO(tie_low_T1Y71));
  sky130_fd_sc_hd__conb_1 conb_T1Y72 (.HI(tie_high_T1Y72), .LO(tie_low_T1Y72));
  sky130_fd_sc_hd__conb_1 conb_T1Y73 (.HI(tie_high_T1Y73), .LO(tie_low_T1Y73));
  sky130_fd_sc_hd__conb_1 conb_T1Y74 (.HI(tie_high_T1Y74), .LO(tie_low_T1Y74));
  sky130_fd_sc_hd__conb_1 conb_T1Y75 (.HI(tie_high_T1Y75), .LO(tie_low_T1Y75));
  sky130_fd_sc_hd__conb_1 conb_T1Y76 (.HI(tie_high_T1Y76), .LO(tie_low_T1Y76));
  sky130_fd_sc_hd__conb_1 conb_T1Y77 (.HI(tie_high_T1Y77), .LO(tie_low_T1Y77));
  sky130_fd_sc_hd__conb_1 conb_T1Y78 (.HI(tie_high_T1Y78), .LO(tie_low_T1Y78));
  sky130_fd_sc_hd__conb_1 conb_T1Y79 (.HI(tie_high_T1Y79), .LO(tie_low_T1Y79));
  sky130_fd_sc_hd__conb_1 conb_T1Y8 (.HI(tie_high_T1Y8), .LO(tie_low_T1Y8));
  sky130_fd_sc_hd__conb_1 conb_T1Y80 (.HI(tie_high_T1Y80), .LO(tie_low_T1Y80));
  sky130_fd_sc_hd__conb_1 conb_T1Y81 (.HI(tie_high_T1Y81), .LO(tie_low_T1Y81));
  sky130_fd_sc_hd__conb_1 conb_T1Y82 (.HI(tie_high_T1Y82), .LO(tie_low_T1Y82));
  sky130_fd_sc_hd__conb_1 conb_T1Y83 (.HI(tie_high_T1Y83), .LO(tie_low_T1Y83));
  sky130_fd_sc_hd__conb_1 conb_T1Y84 (.HI(tie_high_T1Y84), .LO(tie_low_T1Y84));
  sky130_fd_sc_hd__conb_1 conb_T1Y85 (.HI(tie_high_T1Y85), .LO(tie_low_T1Y85));
  sky130_fd_sc_hd__conb_1 conb_T1Y86 (.HI(tie_high_T1Y86), .LO(tie_low_T1Y86));
  sky130_fd_sc_hd__conb_1 conb_T1Y87 (.HI(tie_high_T1Y87), .LO(tie_low_T1Y87));
  sky130_fd_sc_hd__conb_1 conb_T1Y88 (.HI(tie_high_T1Y88), .LO(tie_low_T1Y88));
  sky130_fd_sc_hd__conb_1 conb_T1Y89 (.HI(tie_high_T1Y89), .LO(tie_low_T1Y89));
  sky130_fd_sc_hd__conb_1 conb_T1Y9 (.HI(tie_high_T1Y9), .LO(tie_low_T1Y9));
  sky130_fd_sc_hd__conb_1 conb_T20Y0 (.HI(tie_high_T20Y0), .LO(tie_low_T20Y0));
  sky130_fd_sc_hd__conb_1 conb_T20Y1 (.HI(tie_high_T20Y1), .LO(tie_low_T20Y1));
  sky130_fd_sc_hd__conb_1 conb_T20Y10 (.HI(tie_high_T20Y10), .LO(tie_low_T20Y10));
  sky130_fd_sc_hd__conb_1 conb_T20Y11 (.HI(tie_high_T20Y11), .LO(tie_low_T20Y11));
  sky130_fd_sc_hd__conb_1 conb_T20Y12 (.HI(tie_high_T20Y12), .LO(tie_low_T20Y12));
  sky130_fd_sc_hd__conb_1 conb_T20Y13 (.HI(tie_high_T20Y13), .LO(tie_low_T20Y13));
  sky130_fd_sc_hd__conb_1 conb_T20Y14 (.HI(tie_high_T20Y14), .LO(tie_low_T20Y14));
  sky130_fd_sc_hd__conb_1 conb_T20Y15 (.HI(tie_high_T20Y15), .LO(tie_low_T20Y15));
  sky130_fd_sc_hd__conb_1 conb_T20Y16 (.HI(tie_high_T20Y16), .LO(tie_low_T20Y16));
  sky130_fd_sc_hd__conb_1 conb_T20Y17 (.HI(tie_high_T20Y17), .LO(tie_low_T20Y17));
  sky130_fd_sc_hd__conb_1 conb_T20Y18 (.HI(tie_high_T20Y18), .LO(tie_low_T20Y18));
  sky130_fd_sc_hd__conb_1 conb_T20Y19 (.HI(tie_high_T20Y19), .LO(tie_low_T20Y19));
  sky130_fd_sc_hd__conb_1 conb_T20Y2 (.HI(tie_high_T20Y2), .LO(tie_low_T20Y2));
  sky130_fd_sc_hd__conb_1 conb_T20Y20 (.HI(tie_high_T20Y20), .LO(tie_low_T20Y20));
  sky130_fd_sc_hd__conb_1 conb_T20Y21 (.HI(tie_high_T20Y21), .LO(tie_low_T20Y21));
  sky130_fd_sc_hd__conb_1 conb_T20Y22 (.HI(tie_high_T20Y22), .LO(tie_low_T20Y22));
  sky130_fd_sc_hd__conb_1 conb_T20Y23 (.HI(tie_high_T20Y23), .LO(tie_low_T20Y23));
  sky130_fd_sc_hd__conb_1 conb_T20Y24 (.HI(tie_high_T20Y24), .LO(tie_low_T20Y24));
  sky130_fd_sc_hd__conb_1 conb_T20Y25 (.HI(tie_high_T20Y25), .LO(tie_low_T20Y25));
  sky130_fd_sc_hd__conb_1 conb_T20Y26 (.HI(tie_high_T20Y26), .LO(tie_low_T20Y26));
  sky130_fd_sc_hd__conb_1 conb_T20Y27 (.HI(tie_high_T20Y27), .LO(tie_low_T20Y27));
  sky130_fd_sc_hd__conb_1 conb_T20Y28 (.HI(tie_high_T20Y28), .LO(tie_low_T20Y28));
  sky130_fd_sc_hd__conb_1 conb_T20Y29 (.HI(tie_high_T20Y29), .LO(tie_low_T20Y29));
  sky130_fd_sc_hd__conb_1 conb_T20Y3 (.HI(tie_high_T20Y3), .LO(tie_low_T20Y3));
  sky130_fd_sc_hd__conb_1 conb_T20Y30 (.HI(tie_high_T20Y30), .LO(tie_low_T20Y30));
  sky130_fd_sc_hd__conb_1 conb_T20Y31 (.HI(tie_high_T20Y31), .LO(tie_low_T20Y31));
  sky130_fd_sc_hd__conb_1 conb_T20Y32 (.HI(tie_high_T20Y32), .LO(tie_low_T20Y32));
  sky130_fd_sc_hd__conb_1 conb_T20Y33 (.HI(tie_high_T20Y33), .LO(tie_low_T20Y33));
  sky130_fd_sc_hd__conb_1 conb_T20Y34 (.HI(tie_high_T20Y34), .LO(tie_low_T20Y34));
  sky130_fd_sc_hd__conb_1 conb_T20Y35 (.HI(tie_high_T20Y35), .LO(tie_low_T20Y35));
  sky130_fd_sc_hd__conb_1 conb_T20Y36 (.HI(tie_high_T20Y36), .LO(tie_low_T20Y36));
  sky130_fd_sc_hd__conb_1 conb_T20Y37 (.HI(tie_high_T20Y37), .LO(tie_low_T20Y37));
  sky130_fd_sc_hd__conb_1 conb_T20Y38 (.HI(tie_high_T20Y38), .LO(tie_low_T20Y38));
  sky130_fd_sc_hd__conb_1 conb_T20Y39 (.HI(tie_high_T20Y39), .LO(tie_low_T20Y39));
  sky130_fd_sc_hd__conb_1 conb_T20Y4 (.HI(tie_high_T20Y4), .LO(tie_low_T20Y4));
  sky130_fd_sc_hd__conb_1 conb_T20Y40 (.HI(tie_high_T20Y40), .LO(tie_low_T20Y40));
  sky130_fd_sc_hd__conb_1 conb_T20Y41 (.HI(tie_high_T20Y41), .LO(tie_low_T20Y41));
  sky130_fd_sc_hd__conb_1 conb_T20Y42 (.HI(tie_high_T20Y42), .LO(tie_low_T20Y42));
  sky130_fd_sc_hd__conb_1 conb_T20Y43 (.HI(tie_high_T20Y43), .LO(tie_low_T20Y43));
  sky130_fd_sc_hd__conb_1 conb_T20Y44 (.HI(tie_high_T20Y44), .LO(tie_low_T20Y44));
  sky130_fd_sc_hd__conb_1 conb_T20Y45 (.HI(tie_high_T20Y45), .LO(tie_low_T20Y45));
  sky130_fd_sc_hd__conb_1 conb_T20Y46 (.HI(tie_high_T20Y46), .LO(tie_low_T20Y46));
  sky130_fd_sc_hd__conb_1 conb_T20Y47 (.HI(tie_high_T20Y47), .LO(tie_low_T20Y47));
  sky130_fd_sc_hd__conb_1 conb_T20Y48 (.HI(tie_high_T20Y48), .LO(tie_low_T20Y48));
  sky130_fd_sc_hd__conb_1 conb_T20Y49 (.HI(tie_high_T20Y49), .LO(tie_low_T20Y49));
  sky130_fd_sc_hd__conb_1 conb_T20Y5 (.HI(tie_high_T20Y5), .LO(tie_low_T20Y5));
  sky130_fd_sc_hd__conb_1 conb_T20Y50 (.HI(tie_high_T20Y50), .LO(tie_low_T20Y50));
  sky130_fd_sc_hd__conb_1 conb_T20Y51 (.HI(tie_high_T20Y51), .LO(tie_low_T20Y51));
  sky130_fd_sc_hd__conb_1 conb_T20Y52 (.HI(tie_high_T20Y52), .LO(tie_low_T20Y52));
  sky130_fd_sc_hd__conb_1 conb_T20Y53 (.HI(tie_high_T20Y53), .LO(tie_low_T20Y53));
  sky130_fd_sc_hd__conb_1 conb_T20Y54 (.HI(tie_high_T20Y54), .LO(tie_low_T20Y54));
  sky130_fd_sc_hd__conb_1 conb_T20Y55 (.HI(tie_high_T20Y55), .LO(tie_low_T20Y55));
  sky130_fd_sc_hd__conb_1 conb_T20Y56 (.HI(tie_high_T20Y56), .LO(tie_low_T20Y56));
  sky130_fd_sc_hd__conb_1 conb_T20Y57 (.HI(tie_high_T20Y57), .LO(tie_low_T20Y57));
  sky130_fd_sc_hd__conb_1 conb_T20Y58 (.HI(tie_high_T20Y58), .LO(tie_low_T20Y58));
  sky130_fd_sc_hd__conb_1 conb_T20Y59 (.HI(tie_high_T20Y59), .LO(tie_low_T20Y59));
  sky130_fd_sc_hd__conb_1 conb_T20Y6 (.HI(tie_high_T20Y6), .LO(tie_low_T20Y6));
  sky130_fd_sc_hd__conb_1 conb_T20Y60 (.HI(tie_high_T20Y60), .LO(tie_low_T20Y60));
  sky130_fd_sc_hd__conb_1 conb_T20Y61 (.HI(tie_high_T20Y61), .LO(tie_low_T20Y61));
  sky130_fd_sc_hd__conb_1 conb_T20Y62 (.HI(tie_high_T20Y62), .LO(tie_low_T20Y62));
  sky130_fd_sc_hd__conb_1 conb_T20Y63 (.HI(tie_high_T20Y63), .LO(tie_low_T20Y63));
  sky130_fd_sc_hd__conb_1 conb_T20Y64 (.HI(tie_high_T20Y64), .LO(tie_low_T20Y64));
  sky130_fd_sc_hd__conb_1 conb_T20Y65 (.HI(tie_high_T20Y65), .LO(tie_low_T20Y65));
  sky130_fd_sc_hd__conb_1 conb_T20Y66 (.HI(tie_high_T20Y66), .LO(tie_low_T20Y66));
  sky130_fd_sc_hd__conb_1 conb_T20Y67 (.HI(tie_high_T20Y67), .LO(tie_low_T20Y67));
  sky130_fd_sc_hd__conb_1 conb_T20Y68 (.HI(tie_high_T20Y68), .LO(tie_low_T20Y68));
  sky130_fd_sc_hd__conb_1 conb_T20Y69 (.HI(tie_high_T20Y69), .LO(tie_low_T20Y69));
  sky130_fd_sc_hd__conb_1 conb_T20Y7 (.HI(tie_high_T20Y7), .LO(tie_low_T20Y7));
  sky130_fd_sc_hd__conb_1 conb_T20Y70 (.HI(tie_high_T20Y70), .LO(tie_low_T20Y70));
  sky130_fd_sc_hd__conb_1 conb_T20Y71 (.HI(tie_high_T20Y71), .LO(tie_low_T20Y71));
  sky130_fd_sc_hd__conb_1 conb_T20Y72 (.HI(tie_high_T20Y72), .LO(tie_low_T20Y72));
  sky130_fd_sc_hd__conb_1 conb_T20Y73 (.HI(tie_high_T20Y73), .LO(tie_low_T20Y73));
  sky130_fd_sc_hd__conb_1 conb_T20Y74 (.HI(tie_high_T20Y74), .LO(tie_low_T20Y74));
  sky130_fd_sc_hd__conb_1 conb_T20Y75 (.HI(tie_high_T20Y75), .LO(tie_low_T20Y75));
  sky130_fd_sc_hd__conb_1 conb_T20Y76 (.HI(tie_high_T20Y76), .LO(tie_low_T20Y76));
  sky130_fd_sc_hd__conb_1 conb_T20Y77 (.HI(tie_high_T20Y77), .LO(tie_low_T20Y77));
  sky130_fd_sc_hd__conb_1 conb_T20Y78 (.HI(tie_high_T20Y78), .LO(tie_low_T20Y78));
  sky130_fd_sc_hd__conb_1 conb_T20Y79 (.HI(tie_high_T20Y79), .LO(tie_low_T20Y79));
  sky130_fd_sc_hd__conb_1 conb_T20Y8 (.HI(tie_high_T20Y8), .LO(tie_low_T20Y8));
  sky130_fd_sc_hd__conb_1 conb_T20Y80 (.HI(tie_high_T20Y80), .LO(tie_low_T20Y80));
  sky130_fd_sc_hd__conb_1 conb_T20Y81 (.HI(tie_high_T20Y81), .LO(tie_low_T20Y81));
  sky130_fd_sc_hd__conb_1 conb_T20Y82 (.HI(tie_high_T20Y82), .LO(tie_low_T20Y82));
  sky130_fd_sc_hd__conb_1 conb_T20Y83 (.HI(tie_high_T20Y83), .LO(tie_low_T20Y83));
  sky130_fd_sc_hd__conb_1 conb_T20Y84 (.HI(tie_high_T20Y84), .LO(tie_low_T20Y84));
  sky130_fd_sc_hd__conb_1 conb_T20Y85 (.HI(tie_high_T20Y85), .LO(tie_low_T20Y85));
  sky130_fd_sc_hd__conb_1 conb_T20Y86 (.HI(tie_high_T20Y86), .LO(tie_low_T20Y86));
  sky130_fd_sc_hd__conb_1 conb_T20Y87 (.HI(tie_high_T20Y87), .LO(tie_low_T20Y87));
  sky130_fd_sc_hd__conb_1 conb_T20Y88 (.HI(tie_high_T20Y88), .LO(tie_low_T20Y88));
  sky130_fd_sc_hd__conb_1 conb_T20Y89 (.HI(tie_high_T20Y89), .LO(tie_low_T20Y89));
  sky130_fd_sc_hd__conb_1 conb_T20Y9 (.HI(tie_high_T20Y9), .LO(tie_low_T20Y9));
  sky130_fd_sc_hd__conb_1 conb_T21Y0 (.HI(tie_high_T21Y0), .LO(tie_low_T21Y0));
  sky130_fd_sc_hd__conb_1 conb_T21Y1 (.HI(tie_high_T21Y1), .LO(tie_low_T21Y1));
  sky130_fd_sc_hd__conb_1 conb_T21Y10 (.HI(tie_high_T21Y10), .LO(tie_low_T21Y10));
  sky130_fd_sc_hd__conb_1 conb_T21Y11 (.HI(tie_high_T21Y11), .LO(tie_low_T21Y11));
  sky130_fd_sc_hd__conb_1 conb_T21Y12 (.HI(tie_high_T21Y12), .LO(tie_low_T21Y12));
  sky130_fd_sc_hd__conb_1 conb_T21Y13 (.HI(tie_high_T21Y13), .LO(tie_low_T21Y13));
  sky130_fd_sc_hd__conb_1 conb_T21Y14 (.HI(tie_high_T21Y14), .LO(tie_low_T21Y14));
  sky130_fd_sc_hd__conb_1 conb_T21Y15 (.HI(tie_high_T21Y15), .LO(tie_low_T21Y15));
  sky130_fd_sc_hd__conb_1 conb_T21Y16 (.HI(tie_high_T21Y16), .LO(tie_low_T21Y16));
  sky130_fd_sc_hd__conb_1 conb_T21Y17 (.HI(tie_high_T21Y17), .LO(tie_low_T21Y17));
  sky130_fd_sc_hd__conb_1 conb_T21Y18 (.HI(tie_high_T21Y18), .LO(tie_low_T21Y18));
  sky130_fd_sc_hd__conb_1 conb_T21Y19 (.HI(tie_high_T21Y19), .LO(tie_low_T21Y19));
  sky130_fd_sc_hd__conb_1 conb_T21Y2 (.HI(tie_high_T21Y2), .LO(tie_low_T21Y2));
  sky130_fd_sc_hd__conb_1 conb_T21Y20 (.HI(tie_high_T21Y20), .LO(tie_low_T21Y20));
  sky130_fd_sc_hd__conb_1 conb_T21Y21 (.HI(tie_high_T21Y21), .LO(tie_low_T21Y21));
  sky130_fd_sc_hd__conb_1 conb_T21Y22 (.HI(tie_high_T21Y22), .LO(tie_low_T21Y22));
  sky130_fd_sc_hd__conb_1 conb_T21Y23 (.HI(tie_high_T21Y23), .LO(tie_low_T21Y23));
  sky130_fd_sc_hd__conb_1 conb_T21Y24 (.HI(tie_high_T21Y24), .LO(tie_low_T21Y24));
  sky130_fd_sc_hd__conb_1 conb_T21Y25 (.HI(tie_high_T21Y25), .LO(tie_low_T21Y25));
  sky130_fd_sc_hd__conb_1 conb_T21Y26 (.HI(tie_high_T21Y26), .LO(tie_low_T21Y26));
  sky130_fd_sc_hd__conb_1 conb_T21Y27 (.HI(tie_high_T21Y27), .LO(tie_low_T21Y27));
  sky130_fd_sc_hd__conb_1 conb_T21Y28 (.HI(tie_high_T21Y28), .LO(tie_low_T21Y28));
  sky130_fd_sc_hd__conb_1 conb_T21Y29 (.HI(tie_high_T21Y29), .LO(tie_low_T21Y29));
  sky130_fd_sc_hd__conb_1 conb_T21Y3 (.HI(tie_high_T21Y3), .LO(tie_low_T21Y3));
  sky130_fd_sc_hd__conb_1 conb_T21Y30 (.HI(tie_high_T21Y30), .LO(tie_low_T21Y30));
  sky130_fd_sc_hd__conb_1 conb_T21Y31 (.HI(tie_high_T21Y31), .LO(tie_low_T21Y31));
  sky130_fd_sc_hd__conb_1 conb_T21Y32 (.HI(tie_high_T21Y32), .LO(tie_low_T21Y32));
  sky130_fd_sc_hd__conb_1 conb_T21Y33 (.HI(tie_high_T21Y33), .LO(tie_low_T21Y33));
  sky130_fd_sc_hd__conb_1 conb_T21Y34 (.HI(tie_high_T21Y34), .LO(tie_low_T21Y34));
  sky130_fd_sc_hd__conb_1 conb_T21Y35 (.HI(tie_high_T21Y35), .LO(tie_low_T21Y35));
  sky130_fd_sc_hd__conb_1 conb_T21Y36 (.HI(tie_high_T21Y36), .LO(tie_low_T21Y36));
  sky130_fd_sc_hd__conb_1 conb_T21Y37 (.HI(tie_high_T21Y37), .LO(tie_low_T21Y37));
  sky130_fd_sc_hd__conb_1 conb_T21Y38 (.HI(tie_high_T21Y38), .LO(tie_low_T21Y38));
  sky130_fd_sc_hd__conb_1 conb_T21Y39 (.HI(tie_high_T21Y39), .LO(tie_low_T21Y39));
  sky130_fd_sc_hd__conb_1 conb_T21Y4 (.HI(tie_high_T21Y4), .LO(tie_low_T21Y4));
  sky130_fd_sc_hd__conb_1 conb_T21Y40 (.HI(tie_high_T21Y40), .LO(tie_low_T21Y40));
  sky130_fd_sc_hd__conb_1 conb_T21Y41 (.HI(tie_high_T21Y41), .LO(tie_low_T21Y41));
  sky130_fd_sc_hd__conb_1 conb_T21Y42 (.HI(tie_high_T21Y42), .LO(tie_low_T21Y42));
  sky130_fd_sc_hd__conb_1 conb_T21Y43 (.HI(tie_high_T21Y43), .LO(tie_low_T21Y43));
  sky130_fd_sc_hd__conb_1 conb_T21Y44 (.HI(tie_high_T21Y44), .LO(tie_low_T21Y44));
  sky130_fd_sc_hd__conb_1 conb_T21Y45 (.HI(tie_high_T21Y45), .LO(tie_low_T21Y45));
  sky130_fd_sc_hd__conb_1 conb_T21Y46 (.HI(tie_high_T21Y46), .LO(tie_low_T21Y46));
  sky130_fd_sc_hd__conb_1 conb_T21Y47 (.HI(tie_high_T21Y47), .LO(tie_low_T21Y47));
  sky130_fd_sc_hd__conb_1 conb_T21Y48 (.HI(tie_high_T21Y48), .LO(tie_low_T21Y48));
  sky130_fd_sc_hd__conb_1 conb_T21Y49 (.HI(tie_high_T21Y49), .LO(tie_low_T21Y49));
  sky130_fd_sc_hd__conb_1 conb_T21Y5 (.HI(tie_high_T21Y5), .LO(tie_low_T21Y5));
  sky130_fd_sc_hd__conb_1 conb_T21Y50 (.HI(tie_high_T21Y50), .LO(tie_low_T21Y50));
  sky130_fd_sc_hd__conb_1 conb_T21Y51 (.HI(tie_high_T21Y51), .LO(tie_low_T21Y51));
  sky130_fd_sc_hd__conb_1 conb_T21Y52 (.HI(tie_high_T21Y52), .LO(tie_low_T21Y52));
  sky130_fd_sc_hd__conb_1 conb_T21Y53 (.HI(tie_high_T21Y53), .LO(tie_low_T21Y53));
  sky130_fd_sc_hd__conb_1 conb_T21Y54 (.HI(tie_high_T21Y54), .LO(tie_low_T21Y54));
  sky130_fd_sc_hd__conb_1 conb_T21Y55 (.HI(tie_high_T21Y55), .LO(tie_low_T21Y55));
  sky130_fd_sc_hd__conb_1 conb_T21Y56 (.HI(tie_high_T21Y56), .LO(tie_low_T21Y56));
  sky130_fd_sc_hd__conb_1 conb_T21Y57 (.HI(tie_high_T21Y57), .LO(tie_low_T21Y57));
  sky130_fd_sc_hd__conb_1 conb_T21Y58 (.HI(tie_high_T21Y58), .LO(tie_low_T21Y58));
  sky130_fd_sc_hd__conb_1 conb_T21Y59 (.HI(tie_high_T21Y59), .LO(tie_low_T21Y59));
  sky130_fd_sc_hd__conb_1 conb_T21Y6 (.HI(tie_high_T21Y6), .LO(tie_low_T21Y6));
  sky130_fd_sc_hd__conb_1 conb_T21Y60 (.HI(tie_high_T21Y60), .LO(tie_low_T21Y60));
  sky130_fd_sc_hd__conb_1 conb_T21Y61 (.HI(tie_high_T21Y61), .LO(tie_low_T21Y61));
  sky130_fd_sc_hd__conb_1 conb_T21Y62 (.HI(tie_high_T21Y62), .LO(tie_low_T21Y62));
  sky130_fd_sc_hd__conb_1 conb_T21Y63 (.HI(tie_high_T21Y63), .LO(tie_low_T21Y63));
  sky130_fd_sc_hd__conb_1 conb_T21Y64 (.HI(tie_high_T21Y64), .LO(tie_low_T21Y64));
  sky130_fd_sc_hd__conb_1 conb_T21Y65 (.HI(tie_high_T21Y65), .LO(tie_low_T21Y65));
  sky130_fd_sc_hd__conb_1 conb_T21Y66 (.HI(tie_high_T21Y66), .LO(tie_low_T21Y66));
  sky130_fd_sc_hd__conb_1 conb_T21Y67 (.HI(tie_high_T21Y67), .LO(tie_low_T21Y67));
  sky130_fd_sc_hd__conb_1 conb_T21Y68 (.HI(tie_high_T21Y68), .LO(tie_low_T21Y68));
  sky130_fd_sc_hd__conb_1 conb_T21Y69 (.HI(tie_high_T21Y69), .LO(tie_low_T21Y69));
  sky130_fd_sc_hd__conb_1 conb_T21Y7 (.HI(tie_high_T21Y7), .LO(tie_low_T21Y7));
  sky130_fd_sc_hd__conb_1 conb_T21Y70 (.HI(tie_high_T21Y70), .LO(tie_low_T21Y70));
  sky130_fd_sc_hd__conb_1 conb_T21Y71 (.HI(tie_high_T21Y71), .LO(tie_low_T21Y71));
  sky130_fd_sc_hd__conb_1 conb_T21Y72 (.HI(tie_high_T21Y72), .LO(tie_low_T21Y72));
  sky130_fd_sc_hd__conb_1 conb_T21Y73 (.HI(tie_high_T21Y73), .LO(tie_low_T21Y73));
  sky130_fd_sc_hd__conb_1 conb_T21Y74 (.HI(tie_high_T21Y74), .LO(tie_low_T21Y74));
  sky130_fd_sc_hd__conb_1 conb_T21Y75 (.HI(tie_high_T21Y75), .LO(tie_low_T21Y75));
  sky130_fd_sc_hd__conb_1 conb_T21Y76 (.HI(tie_high_T21Y76), .LO(tie_low_T21Y76));
  sky130_fd_sc_hd__conb_1 conb_T21Y77 (.HI(tie_high_T21Y77), .LO(tie_low_T21Y77));
  sky130_fd_sc_hd__conb_1 conb_T21Y78 (.HI(tie_high_T21Y78), .LO(tie_low_T21Y78));
  sky130_fd_sc_hd__conb_1 conb_T21Y79 (.HI(tie_high_T21Y79), .LO(tie_low_T21Y79));
  sky130_fd_sc_hd__conb_1 conb_T21Y8 (.HI(tie_high_T21Y8), .LO(tie_low_T21Y8));
  sky130_fd_sc_hd__conb_1 conb_T21Y80 (.HI(tie_high_T21Y80), .LO(tie_low_T21Y80));
  sky130_fd_sc_hd__conb_1 conb_T21Y81 (.HI(tie_high_T21Y81), .LO(tie_low_T21Y81));
  sky130_fd_sc_hd__conb_1 conb_T21Y82 (.HI(tie_high_T21Y82), .LO(tie_low_T21Y82));
  sky130_fd_sc_hd__conb_1 conb_T21Y83 (.HI(tie_high_T21Y83), .LO(tie_low_T21Y83));
  sky130_fd_sc_hd__conb_1 conb_T21Y84 (.HI(tie_high_T21Y84), .LO(tie_low_T21Y84));
  sky130_fd_sc_hd__conb_1 conb_T21Y85 (.HI(tie_high_T21Y85), .LO(tie_low_T21Y85));
  sky130_fd_sc_hd__conb_1 conb_T21Y86 (.HI(tie_high_T21Y86), .LO(tie_low_T21Y86));
  sky130_fd_sc_hd__conb_1 conb_T21Y87 (.HI(tie_high_T21Y87), .LO(tie_low_T21Y87));
  sky130_fd_sc_hd__conb_1 conb_T21Y88 (.HI(tie_high_T21Y88), .LO(tie_low_T21Y88));
  sky130_fd_sc_hd__conb_1 conb_T21Y89 (.HI(tie_high_T21Y89), .LO(tie_low_T21Y89));
  sky130_fd_sc_hd__conb_1 conb_T21Y9 (.HI(tie_high_T21Y9), .LO(tie_low_T21Y9));
  sky130_fd_sc_hd__conb_1 conb_T22Y0 (.HI(tie_high_T22Y0), .LO(tie_low_T22Y0));
  sky130_fd_sc_hd__conb_1 conb_T22Y1 (.HI(tie_high_T22Y1), .LO(tie_low_T22Y1));
  sky130_fd_sc_hd__conb_1 conb_T22Y10 (.HI(tie_high_T22Y10), .LO(tie_low_T22Y10));
  sky130_fd_sc_hd__conb_1 conb_T22Y11 (.HI(tie_high_T22Y11), .LO(tie_low_T22Y11));
  sky130_fd_sc_hd__conb_1 conb_T22Y12 (.HI(tie_high_T22Y12), .LO(tie_low_T22Y12));
  sky130_fd_sc_hd__conb_1 conb_T22Y13 (.HI(tie_high_T22Y13), .LO(tie_low_T22Y13));
  sky130_fd_sc_hd__conb_1 conb_T22Y14 (.HI(tie_high_T22Y14), .LO(tie_low_T22Y14));
  sky130_fd_sc_hd__conb_1 conb_T22Y15 (.HI(tie_high_T22Y15), .LO(tie_low_T22Y15));
  sky130_fd_sc_hd__conb_1 conb_T22Y16 (.HI(tie_high_T22Y16), .LO(tie_low_T22Y16));
  sky130_fd_sc_hd__conb_1 conb_T22Y17 (.HI(tie_high_T22Y17), .LO(tie_low_T22Y17));
  sky130_fd_sc_hd__conb_1 conb_T22Y18 (.HI(tie_high_T22Y18), .LO(tie_low_T22Y18));
  sky130_fd_sc_hd__conb_1 conb_T22Y19 (.HI(tie_high_T22Y19), .LO(tie_low_T22Y19));
  sky130_fd_sc_hd__conb_1 conb_T22Y2 (.HI(tie_high_T22Y2), .LO(tie_low_T22Y2));
  sky130_fd_sc_hd__conb_1 conb_T22Y20 (.HI(tie_high_T22Y20), .LO(tie_low_T22Y20));
  sky130_fd_sc_hd__conb_1 conb_T22Y21 (.HI(tie_high_T22Y21), .LO(tie_low_T22Y21));
  sky130_fd_sc_hd__conb_1 conb_T22Y22 (.HI(tie_high_T22Y22), .LO(tie_low_T22Y22));
  sky130_fd_sc_hd__conb_1 conb_T22Y23 (.HI(tie_high_T22Y23), .LO(tie_low_T22Y23));
  sky130_fd_sc_hd__conb_1 conb_T22Y24 (.HI(tie_high_T22Y24), .LO(tie_low_T22Y24));
  sky130_fd_sc_hd__conb_1 conb_T22Y25 (.HI(tie_high_T22Y25), .LO(tie_low_T22Y25));
  sky130_fd_sc_hd__conb_1 conb_T22Y26 (.HI(tie_high_T22Y26), .LO(tie_low_T22Y26));
  sky130_fd_sc_hd__conb_1 conb_T22Y27 (.HI(tie_high_T22Y27), .LO(tie_low_T22Y27));
  sky130_fd_sc_hd__conb_1 conb_T22Y28 (.HI(tie_high_T22Y28), .LO(tie_low_T22Y28));
  sky130_fd_sc_hd__conb_1 conb_T22Y29 (.HI(tie_high_T22Y29), .LO(tie_low_T22Y29));
  sky130_fd_sc_hd__conb_1 conb_T22Y3 (.HI(tie_high_T22Y3), .LO(tie_low_T22Y3));
  sky130_fd_sc_hd__conb_1 conb_T22Y30 (.HI(tie_high_T22Y30), .LO(tie_low_T22Y30));
  sky130_fd_sc_hd__conb_1 conb_T22Y31 (.HI(tie_high_T22Y31), .LO(tie_low_T22Y31));
  sky130_fd_sc_hd__conb_1 conb_T22Y32 (.HI(tie_high_T22Y32), .LO(tie_low_T22Y32));
  sky130_fd_sc_hd__conb_1 conb_T22Y33 (.HI(tie_high_T22Y33), .LO(tie_low_T22Y33));
  sky130_fd_sc_hd__conb_1 conb_T22Y34 (.HI(tie_high_T22Y34), .LO(tie_low_T22Y34));
  sky130_fd_sc_hd__conb_1 conb_T22Y35 (.HI(tie_high_T22Y35), .LO(tie_low_T22Y35));
  sky130_fd_sc_hd__conb_1 conb_T22Y36 (.HI(tie_high_T22Y36), .LO(tie_low_T22Y36));
  sky130_fd_sc_hd__conb_1 conb_T22Y37 (.HI(tie_high_T22Y37), .LO(tie_low_T22Y37));
  sky130_fd_sc_hd__conb_1 conb_T22Y38 (.HI(tie_high_T22Y38), .LO(tie_low_T22Y38));
  sky130_fd_sc_hd__conb_1 conb_T22Y39 (.HI(tie_high_T22Y39), .LO(tie_low_T22Y39));
  sky130_fd_sc_hd__conb_1 conb_T22Y4 (.HI(tie_high_T22Y4), .LO(tie_low_T22Y4));
  sky130_fd_sc_hd__conb_1 conb_T22Y40 (.HI(tie_high_T22Y40), .LO(tie_low_T22Y40));
  sky130_fd_sc_hd__conb_1 conb_T22Y41 (.HI(tie_high_T22Y41), .LO(tie_low_T22Y41));
  sky130_fd_sc_hd__conb_1 conb_T22Y42 (.HI(tie_high_T22Y42), .LO(tie_low_T22Y42));
  sky130_fd_sc_hd__conb_1 conb_T22Y43 (.HI(tie_high_T22Y43), .LO(tie_low_T22Y43));
  sky130_fd_sc_hd__conb_1 conb_T22Y44 (.HI(tie_high_T22Y44), .LO(tie_low_T22Y44));
  sky130_fd_sc_hd__conb_1 conb_T22Y45 (.HI(tie_high_T22Y45), .LO(tie_low_T22Y45));
  sky130_fd_sc_hd__conb_1 conb_T22Y46 (.HI(tie_high_T22Y46), .LO(tie_low_T22Y46));
  sky130_fd_sc_hd__conb_1 conb_T22Y47 (.HI(tie_high_T22Y47), .LO(tie_low_T22Y47));
  sky130_fd_sc_hd__conb_1 conb_T22Y48 (.HI(tie_high_T22Y48), .LO(tie_low_T22Y48));
  sky130_fd_sc_hd__conb_1 conb_T22Y49 (.HI(tie_high_T22Y49), .LO(tie_low_T22Y49));
  sky130_fd_sc_hd__conb_1 conb_T22Y5 (.HI(tie_high_T22Y5), .LO(tie_low_T22Y5));
  sky130_fd_sc_hd__conb_1 conb_T22Y50 (.HI(tie_high_T22Y50), .LO(tie_low_T22Y50));
  sky130_fd_sc_hd__conb_1 conb_T22Y51 (.HI(tie_high_T22Y51), .LO(tie_low_T22Y51));
  sky130_fd_sc_hd__conb_1 conb_T22Y52 (.HI(tie_high_T22Y52), .LO(tie_low_T22Y52));
  sky130_fd_sc_hd__conb_1 conb_T22Y53 (.HI(tie_high_T22Y53), .LO(tie_low_T22Y53));
  sky130_fd_sc_hd__conb_1 conb_T22Y54 (.HI(tie_high_T22Y54), .LO(tie_low_T22Y54));
  sky130_fd_sc_hd__conb_1 conb_T22Y55 (.HI(tie_high_T22Y55), .LO(tie_low_T22Y55));
  sky130_fd_sc_hd__conb_1 conb_T22Y56 (.HI(tie_high_T22Y56), .LO(tie_low_T22Y56));
  sky130_fd_sc_hd__conb_1 conb_T22Y57 (.HI(tie_high_T22Y57), .LO(tie_low_T22Y57));
  sky130_fd_sc_hd__conb_1 conb_T22Y58 (.HI(tie_high_T22Y58), .LO(tie_low_T22Y58));
  sky130_fd_sc_hd__conb_1 conb_T22Y59 (.HI(tie_high_T22Y59), .LO(tie_low_T22Y59));
  sky130_fd_sc_hd__conb_1 conb_T22Y6 (.HI(tie_high_T22Y6), .LO(tie_low_T22Y6));
  sky130_fd_sc_hd__conb_1 conb_T22Y60 (.HI(tie_high_T22Y60), .LO(tie_low_T22Y60));
  sky130_fd_sc_hd__conb_1 conb_T22Y61 (.HI(tie_high_T22Y61), .LO(tie_low_T22Y61));
  sky130_fd_sc_hd__conb_1 conb_T22Y62 (.HI(tie_high_T22Y62), .LO(tie_low_T22Y62));
  sky130_fd_sc_hd__conb_1 conb_T22Y63 (.HI(tie_high_T22Y63), .LO(tie_low_T22Y63));
  sky130_fd_sc_hd__conb_1 conb_T22Y64 (.HI(tie_high_T22Y64), .LO(tie_low_T22Y64));
  sky130_fd_sc_hd__conb_1 conb_T22Y65 (.HI(tie_high_T22Y65), .LO(tie_low_T22Y65));
  sky130_fd_sc_hd__conb_1 conb_T22Y66 (.HI(tie_high_T22Y66), .LO(tie_low_T22Y66));
  sky130_fd_sc_hd__conb_1 conb_T22Y67 (.HI(tie_high_T22Y67), .LO(tie_low_T22Y67));
  sky130_fd_sc_hd__conb_1 conb_T22Y68 (.HI(tie_high_T22Y68), .LO(tie_low_T22Y68));
  sky130_fd_sc_hd__conb_1 conb_T22Y69 (.HI(tie_high_T22Y69), .LO(tie_low_T22Y69));
  sky130_fd_sc_hd__conb_1 conb_T22Y7 (.HI(tie_high_T22Y7), .LO(tie_low_T22Y7));
  sky130_fd_sc_hd__conb_1 conb_T22Y70 (.HI(tie_high_T22Y70), .LO(tie_low_T22Y70));
  sky130_fd_sc_hd__conb_1 conb_T22Y71 (.HI(tie_high_T22Y71), .LO(tie_low_T22Y71));
  sky130_fd_sc_hd__conb_1 conb_T22Y72 (.HI(tie_high_T22Y72), .LO(tie_low_T22Y72));
  sky130_fd_sc_hd__conb_1 conb_T22Y73 (.HI(tie_high_T22Y73), .LO(tie_low_T22Y73));
  sky130_fd_sc_hd__conb_1 conb_T22Y74 (.HI(tie_high_T22Y74), .LO(tie_low_T22Y74));
  sky130_fd_sc_hd__conb_1 conb_T22Y75 (.HI(tie_high_T22Y75), .LO(tie_low_T22Y75));
  sky130_fd_sc_hd__conb_1 conb_T22Y76 (.HI(tie_high_T22Y76), .LO(tie_low_T22Y76));
  sky130_fd_sc_hd__conb_1 conb_T22Y77 (.HI(tie_high_T22Y77), .LO(tie_low_T22Y77));
  sky130_fd_sc_hd__conb_1 conb_T22Y78 (.HI(tie_high_T22Y78), .LO(tie_low_T22Y78));
  sky130_fd_sc_hd__conb_1 conb_T22Y79 (.HI(tie_high_T22Y79), .LO(tie_low_T22Y79));
  sky130_fd_sc_hd__conb_1 conb_T22Y8 (.HI(tie_high_T22Y8), .LO(tie_low_T22Y8));
  sky130_fd_sc_hd__conb_1 conb_T22Y80 (.HI(tie_high_T22Y80), .LO(tie_low_T22Y80));
  sky130_fd_sc_hd__conb_1 conb_T22Y81 (.HI(tie_high_T22Y81), .LO(tie_low_T22Y81));
  sky130_fd_sc_hd__conb_1 conb_T22Y82 (.HI(tie_high_T22Y82), .LO(tie_low_T22Y82));
  sky130_fd_sc_hd__conb_1 conb_T22Y83 (.HI(tie_high_T22Y83), .LO(tie_low_T22Y83));
  sky130_fd_sc_hd__conb_1 conb_T22Y84 (.HI(tie_high_T22Y84), .LO(tie_low_T22Y84));
  sky130_fd_sc_hd__conb_1 conb_T22Y85 (.HI(tie_high_T22Y85), .LO(tie_low_T22Y85));
  sky130_fd_sc_hd__conb_1 conb_T22Y86 (.HI(tie_high_T22Y86), .LO(tie_low_T22Y86));
  sky130_fd_sc_hd__conb_1 conb_T22Y87 (.HI(tie_high_T22Y87), .LO(tie_low_T22Y87));
  sky130_fd_sc_hd__conb_1 conb_T22Y88 (.HI(tie_high_T22Y88), .LO(tie_low_T22Y88));
  sky130_fd_sc_hd__conb_1 conb_T22Y89 (.HI(tie_high_T22Y89), .LO(tie_low_T22Y89));
  sky130_fd_sc_hd__conb_1 conb_T22Y9 (.HI(tie_high_T22Y9), .LO(tie_low_T22Y9));
  sky130_fd_sc_hd__conb_1 conb_T23Y0 (.HI(tie_high_T23Y0), .LO(tie_low_T23Y0));
  sky130_fd_sc_hd__conb_1 conb_T23Y1 (.HI(tie_high_T23Y1), .LO(tie_low_T23Y1));
  sky130_fd_sc_hd__conb_1 conb_T23Y10 (.HI(tie_high_T23Y10), .LO(tie_low_T23Y10));
  sky130_fd_sc_hd__conb_1 conb_T23Y11 (.HI(tie_high_T23Y11), .LO(tie_low_T23Y11));
  sky130_fd_sc_hd__conb_1 conb_T23Y12 (.HI(tie_high_T23Y12), .LO(tie_low_T23Y12));
  sky130_fd_sc_hd__conb_1 conb_T23Y13 (.HI(tie_high_T23Y13), .LO(tie_low_T23Y13));
  sky130_fd_sc_hd__conb_1 conb_T23Y14 (.HI(tie_high_T23Y14), .LO(tie_low_T23Y14));
  sky130_fd_sc_hd__conb_1 conb_T23Y15 (.HI(tie_high_T23Y15), .LO(tie_low_T23Y15));
  sky130_fd_sc_hd__conb_1 conb_T23Y16 (.HI(tie_high_T23Y16), .LO(tie_low_T23Y16));
  sky130_fd_sc_hd__conb_1 conb_T23Y17 (.HI(tie_high_T23Y17), .LO(tie_low_T23Y17));
  sky130_fd_sc_hd__conb_1 conb_T23Y18 (.HI(tie_high_T23Y18), .LO(tie_low_T23Y18));
  sky130_fd_sc_hd__conb_1 conb_T23Y19 (.HI(tie_high_T23Y19), .LO(tie_low_T23Y19));
  sky130_fd_sc_hd__conb_1 conb_T23Y2 (.HI(tie_high_T23Y2), .LO(tie_low_T23Y2));
  sky130_fd_sc_hd__conb_1 conb_T23Y20 (.HI(tie_high_T23Y20), .LO(tie_low_T23Y20));
  sky130_fd_sc_hd__conb_1 conb_T23Y21 (.HI(tie_high_T23Y21), .LO(tie_low_T23Y21));
  sky130_fd_sc_hd__conb_1 conb_T23Y22 (.HI(tie_high_T23Y22), .LO(tie_low_T23Y22));
  sky130_fd_sc_hd__conb_1 conb_T23Y23 (.HI(tie_high_T23Y23), .LO(tie_low_T23Y23));
  sky130_fd_sc_hd__conb_1 conb_T23Y24 (.HI(tie_high_T23Y24), .LO(tie_low_T23Y24));
  sky130_fd_sc_hd__conb_1 conb_T23Y25 (.HI(tie_high_T23Y25), .LO(tie_low_T23Y25));
  sky130_fd_sc_hd__conb_1 conb_T23Y26 (.HI(tie_high_T23Y26), .LO(tie_low_T23Y26));
  sky130_fd_sc_hd__conb_1 conb_T23Y27 (.HI(tie_high_T23Y27), .LO(tie_low_T23Y27));
  sky130_fd_sc_hd__conb_1 conb_T23Y28 (.HI(tie_high_T23Y28), .LO(tie_low_T23Y28));
  sky130_fd_sc_hd__conb_1 conb_T23Y29 (.HI(tie_high_T23Y29), .LO(tie_low_T23Y29));
  sky130_fd_sc_hd__conb_1 conb_T23Y3 (.HI(tie_high_T23Y3), .LO(tie_low_T23Y3));
  sky130_fd_sc_hd__conb_1 conb_T23Y30 (.HI(tie_high_T23Y30), .LO(tie_low_T23Y30));
  sky130_fd_sc_hd__conb_1 conb_T23Y31 (.HI(tie_high_T23Y31), .LO(tie_low_T23Y31));
  sky130_fd_sc_hd__conb_1 conb_T23Y32 (.HI(tie_high_T23Y32), .LO(tie_low_T23Y32));
  sky130_fd_sc_hd__conb_1 conb_T23Y33 (.HI(tie_high_T23Y33), .LO(tie_low_T23Y33));
  sky130_fd_sc_hd__conb_1 conb_T23Y34 (.HI(tie_high_T23Y34), .LO(tie_low_T23Y34));
  sky130_fd_sc_hd__conb_1 conb_T23Y35 (.HI(tie_high_T23Y35), .LO(tie_low_T23Y35));
  sky130_fd_sc_hd__conb_1 conb_T23Y36 (.HI(tie_high_T23Y36), .LO(tie_low_T23Y36));
  sky130_fd_sc_hd__conb_1 conb_T23Y37 (.HI(tie_high_T23Y37), .LO(tie_low_T23Y37));
  sky130_fd_sc_hd__conb_1 conb_T23Y38 (.HI(tie_high_T23Y38), .LO(tie_low_T23Y38));
  sky130_fd_sc_hd__conb_1 conb_T23Y39 (.HI(tie_high_T23Y39), .LO(tie_low_T23Y39));
  sky130_fd_sc_hd__conb_1 conb_T23Y4 (.HI(tie_high_T23Y4), .LO(tie_low_T23Y4));
  sky130_fd_sc_hd__conb_1 conb_T23Y40 (.HI(tie_high_T23Y40), .LO(tie_low_T23Y40));
  sky130_fd_sc_hd__conb_1 conb_T23Y41 (.HI(tie_high_T23Y41), .LO(tie_low_T23Y41));
  sky130_fd_sc_hd__conb_1 conb_T23Y42 (.HI(tie_high_T23Y42), .LO(tie_low_T23Y42));
  sky130_fd_sc_hd__conb_1 conb_T23Y43 (.HI(tie_high_T23Y43), .LO(tie_low_T23Y43));
  sky130_fd_sc_hd__conb_1 conb_T23Y44 (.HI(tie_high_T23Y44), .LO(tie_low_T23Y44));
  sky130_fd_sc_hd__conb_1 conb_T23Y45 (.HI(tie_high_T23Y45), .LO(tie_low_T23Y45));
  sky130_fd_sc_hd__conb_1 conb_T23Y46 (.HI(tie_high_T23Y46), .LO(tie_low_T23Y46));
  sky130_fd_sc_hd__conb_1 conb_T23Y47 (.HI(tie_high_T23Y47), .LO(tie_low_T23Y47));
  sky130_fd_sc_hd__conb_1 conb_T23Y48 (.HI(tie_high_T23Y48), .LO(tie_low_T23Y48));
  sky130_fd_sc_hd__conb_1 conb_T23Y49 (.HI(tie_high_T23Y49), .LO(tie_low_T23Y49));
  sky130_fd_sc_hd__conb_1 conb_T23Y5 (.HI(tie_high_T23Y5), .LO(tie_low_T23Y5));
  sky130_fd_sc_hd__conb_1 conb_T23Y50 (.HI(tie_high_T23Y50), .LO(tie_low_T23Y50));
  sky130_fd_sc_hd__conb_1 conb_T23Y51 (.HI(tie_high_T23Y51), .LO(tie_low_T23Y51));
  sky130_fd_sc_hd__conb_1 conb_T23Y52 (.HI(tie_high_T23Y52), .LO(tie_low_T23Y52));
  sky130_fd_sc_hd__conb_1 conb_T23Y53 (.HI(tie_high_T23Y53), .LO(tie_low_T23Y53));
  sky130_fd_sc_hd__conb_1 conb_T23Y54 (.HI(tie_high_T23Y54), .LO(tie_low_T23Y54));
  sky130_fd_sc_hd__conb_1 conb_T23Y55 (.HI(tie_high_T23Y55), .LO(tie_low_T23Y55));
  sky130_fd_sc_hd__conb_1 conb_T23Y56 (.HI(tie_high_T23Y56), .LO(tie_low_T23Y56));
  sky130_fd_sc_hd__conb_1 conb_T23Y57 (.HI(tie_high_T23Y57), .LO(tie_low_T23Y57));
  sky130_fd_sc_hd__conb_1 conb_T23Y58 (.HI(tie_high_T23Y58), .LO(tie_low_T23Y58));
  sky130_fd_sc_hd__conb_1 conb_T23Y59 (.HI(tie_high_T23Y59), .LO(tie_low_T23Y59));
  sky130_fd_sc_hd__conb_1 conb_T23Y6 (.HI(tie_high_T23Y6), .LO(tie_low_T23Y6));
  sky130_fd_sc_hd__conb_1 conb_T23Y60 (.HI(tie_high_T23Y60), .LO(tie_low_T23Y60));
  sky130_fd_sc_hd__conb_1 conb_T23Y61 (.HI(tie_high_T23Y61), .LO(tie_low_T23Y61));
  sky130_fd_sc_hd__conb_1 conb_T23Y62 (.HI(tie_high_T23Y62), .LO(tie_low_T23Y62));
  sky130_fd_sc_hd__conb_1 conb_T23Y63 (.HI(tie_high_T23Y63), .LO(tie_low_T23Y63));
  sky130_fd_sc_hd__conb_1 conb_T23Y64 (.HI(tie_high_T23Y64), .LO(tie_low_T23Y64));
  sky130_fd_sc_hd__conb_1 conb_T23Y65 (.HI(tie_high_T23Y65), .LO(tie_low_T23Y65));
  sky130_fd_sc_hd__conb_1 conb_T23Y66 (.HI(tie_high_T23Y66), .LO(tie_low_T23Y66));
  sky130_fd_sc_hd__conb_1 conb_T23Y67 (.HI(tie_high_T23Y67), .LO(tie_low_T23Y67));
  sky130_fd_sc_hd__conb_1 conb_T23Y68 (.HI(tie_high_T23Y68), .LO(tie_low_T23Y68));
  sky130_fd_sc_hd__conb_1 conb_T23Y69 (.HI(tie_high_T23Y69), .LO(tie_low_T23Y69));
  sky130_fd_sc_hd__conb_1 conb_T23Y7 (.HI(tie_high_T23Y7), .LO(tie_low_T23Y7));
  sky130_fd_sc_hd__conb_1 conb_T23Y70 (.HI(tie_high_T23Y70), .LO(tie_low_T23Y70));
  sky130_fd_sc_hd__conb_1 conb_T23Y71 (.HI(tie_high_T23Y71), .LO(tie_low_T23Y71));
  sky130_fd_sc_hd__conb_1 conb_T23Y72 (.HI(tie_high_T23Y72), .LO(tie_low_T23Y72));
  sky130_fd_sc_hd__conb_1 conb_T23Y73 (.HI(tie_high_T23Y73), .LO(tie_low_T23Y73));
  sky130_fd_sc_hd__conb_1 conb_T23Y74 (.HI(tie_high_T23Y74), .LO(tie_low_T23Y74));
  sky130_fd_sc_hd__conb_1 conb_T23Y75 (.HI(tie_high_T23Y75), .LO(tie_low_T23Y75));
  sky130_fd_sc_hd__conb_1 conb_T23Y76 (.HI(tie_high_T23Y76), .LO(tie_low_T23Y76));
  sky130_fd_sc_hd__conb_1 conb_T23Y77 (.HI(tie_high_T23Y77), .LO(tie_low_T23Y77));
  sky130_fd_sc_hd__conb_1 conb_T23Y78 (.HI(tie_high_T23Y78), .LO(tie_low_T23Y78));
  sky130_fd_sc_hd__conb_1 conb_T23Y79 (.HI(tie_high_T23Y79), .LO(tie_low_T23Y79));
  sky130_fd_sc_hd__conb_1 conb_T23Y8 (.HI(tie_high_T23Y8), .LO(tie_low_T23Y8));
  sky130_fd_sc_hd__conb_1 conb_T23Y80 (.HI(tie_high_T23Y80), .LO(tie_low_T23Y80));
  sky130_fd_sc_hd__conb_1 conb_T23Y81 (.HI(tie_high_T23Y81), .LO(tie_low_T23Y81));
  sky130_fd_sc_hd__conb_1 conb_T23Y82 (.HI(tie_high_T23Y82), .LO(tie_low_T23Y82));
  sky130_fd_sc_hd__conb_1 conb_T23Y83 (.HI(tie_high_T23Y83), .LO(tie_low_T23Y83));
  sky130_fd_sc_hd__conb_1 conb_T23Y84 (.HI(tie_high_T23Y84), .LO(tie_low_T23Y84));
  sky130_fd_sc_hd__conb_1 conb_T23Y85 (.HI(tie_high_T23Y85), .LO(tie_low_T23Y85));
  sky130_fd_sc_hd__conb_1 conb_T23Y86 (.HI(tie_high_T23Y86), .LO(tie_low_T23Y86));
  sky130_fd_sc_hd__conb_1 conb_T23Y87 (.HI(tie_high_T23Y87), .LO(tie_low_T23Y87));
  sky130_fd_sc_hd__conb_1 conb_T23Y88 (.HI(tie_high_T23Y88), .LO(tie_low_T23Y88));
  sky130_fd_sc_hd__conb_1 conb_T23Y89 (.HI(tie_high_T23Y89), .LO(tie_low_T23Y89));
  sky130_fd_sc_hd__conb_1 conb_T23Y9 (.HI(tie_high_T23Y9), .LO(tie_low_T23Y9));
  sky130_fd_sc_hd__conb_1 conb_T24Y0 (.HI(tie_high_T24Y0), .LO(tie_low_T24Y0));
  sky130_fd_sc_hd__conb_1 conb_T24Y1 (.HI(tie_high_T24Y1), .LO(tie_low_T24Y1));
  sky130_fd_sc_hd__conb_1 conb_T24Y10 (.HI(tie_high_T24Y10), .LO(tie_low_T24Y10));
  sky130_fd_sc_hd__conb_1 conb_T24Y11 (.HI(tie_high_T24Y11), .LO(tie_low_T24Y11));
  sky130_fd_sc_hd__conb_1 conb_T24Y12 (.HI(tie_high_T24Y12), .LO(tie_low_T24Y12));
  sky130_fd_sc_hd__conb_1 conb_T24Y13 (.HI(tie_high_T24Y13), .LO(tie_low_T24Y13));
  sky130_fd_sc_hd__conb_1 conb_T24Y14 (.HI(tie_high_T24Y14), .LO(tie_low_T24Y14));
  sky130_fd_sc_hd__conb_1 conb_T24Y15 (.HI(tie_high_T24Y15), .LO(tie_low_T24Y15));
  sky130_fd_sc_hd__conb_1 conb_T24Y16 (.HI(tie_high_T24Y16), .LO(tie_low_T24Y16));
  sky130_fd_sc_hd__conb_1 conb_T24Y17 (.HI(tie_high_T24Y17), .LO(tie_low_T24Y17));
  sky130_fd_sc_hd__conb_1 conb_T24Y18 (.HI(tie_high_T24Y18), .LO(tie_low_T24Y18));
  sky130_fd_sc_hd__conb_1 conb_T24Y19 (.HI(tie_high_T24Y19), .LO(tie_low_T24Y19));
  sky130_fd_sc_hd__conb_1 conb_T24Y2 (.HI(tie_high_T24Y2), .LO(tie_low_T24Y2));
  sky130_fd_sc_hd__conb_1 conb_T24Y20 (.HI(tie_high_T24Y20), .LO(tie_low_T24Y20));
  sky130_fd_sc_hd__conb_1 conb_T24Y21 (.HI(tie_high_T24Y21), .LO(tie_low_T24Y21));
  sky130_fd_sc_hd__conb_1 conb_T24Y22 (.HI(tie_high_T24Y22), .LO(tie_low_T24Y22));
  sky130_fd_sc_hd__conb_1 conb_T24Y23 (.HI(tie_high_T24Y23), .LO(tie_low_T24Y23));
  sky130_fd_sc_hd__conb_1 conb_T24Y24 (.HI(tie_high_T24Y24), .LO(tie_low_T24Y24));
  sky130_fd_sc_hd__conb_1 conb_T24Y25 (.HI(tie_high_T24Y25), .LO(tie_low_T24Y25));
  sky130_fd_sc_hd__conb_1 conb_T24Y26 (.HI(tie_high_T24Y26), .LO(tie_low_T24Y26));
  sky130_fd_sc_hd__conb_1 conb_T24Y27 (.HI(tie_high_T24Y27), .LO(tie_low_T24Y27));
  sky130_fd_sc_hd__conb_1 conb_T24Y28 (.HI(tie_high_T24Y28), .LO(tie_low_T24Y28));
  sky130_fd_sc_hd__conb_1 conb_T24Y29 (.HI(tie_high_T24Y29), .LO(tie_low_T24Y29));
  sky130_fd_sc_hd__conb_1 conb_T24Y3 (.HI(tie_high_T24Y3), .LO(tie_low_T24Y3));
  sky130_fd_sc_hd__conb_1 conb_T24Y30 (.HI(tie_high_T24Y30), .LO(tie_low_T24Y30));
  sky130_fd_sc_hd__conb_1 conb_T24Y31 (.HI(tie_high_T24Y31), .LO(tie_low_T24Y31));
  sky130_fd_sc_hd__conb_1 conb_T24Y32 (.HI(tie_high_T24Y32), .LO(tie_low_T24Y32));
  sky130_fd_sc_hd__conb_1 conb_T24Y33 (.HI(tie_high_T24Y33), .LO(tie_low_T24Y33));
  sky130_fd_sc_hd__conb_1 conb_T24Y34 (.HI(tie_high_T24Y34), .LO(tie_low_T24Y34));
  sky130_fd_sc_hd__conb_1 conb_T24Y35 (.HI(tie_high_T24Y35), .LO(tie_low_T24Y35));
  sky130_fd_sc_hd__conb_1 conb_T24Y36 (.HI(tie_high_T24Y36), .LO(tie_low_T24Y36));
  sky130_fd_sc_hd__conb_1 conb_T24Y37 (.HI(tie_high_T24Y37), .LO(tie_low_T24Y37));
  sky130_fd_sc_hd__conb_1 conb_T24Y38 (.HI(tie_high_T24Y38), .LO(tie_low_T24Y38));
  sky130_fd_sc_hd__conb_1 conb_T24Y39 (.HI(tie_high_T24Y39), .LO(tie_low_T24Y39));
  sky130_fd_sc_hd__conb_1 conb_T24Y4 (.HI(tie_high_T24Y4), .LO(tie_low_T24Y4));
  sky130_fd_sc_hd__conb_1 conb_T24Y40 (.HI(tie_high_T24Y40), .LO(tie_low_T24Y40));
  sky130_fd_sc_hd__conb_1 conb_T24Y41 (.HI(tie_high_T24Y41), .LO(tie_low_T24Y41));
  sky130_fd_sc_hd__conb_1 conb_T24Y42 (.HI(tie_high_T24Y42), .LO(tie_low_T24Y42));
  sky130_fd_sc_hd__conb_1 conb_T24Y43 (.HI(tie_high_T24Y43), .LO(tie_low_T24Y43));
  sky130_fd_sc_hd__conb_1 conb_T24Y44 (.HI(tie_high_T24Y44), .LO(tie_low_T24Y44));
  sky130_fd_sc_hd__conb_1 conb_T24Y45 (.HI(tie_high_T24Y45), .LO(tie_low_T24Y45));
  sky130_fd_sc_hd__conb_1 conb_T24Y46 (.HI(tie_high_T24Y46), .LO(tie_low_T24Y46));
  sky130_fd_sc_hd__conb_1 conb_T24Y47 (.HI(tie_high_T24Y47), .LO(tie_low_T24Y47));
  sky130_fd_sc_hd__conb_1 conb_T24Y48 (.HI(tie_high_T24Y48), .LO(tie_low_T24Y48));
  sky130_fd_sc_hd__conb_1 conb_T24Y49 (.HI(tie_high_T24Y49), .LO(tie_low_T24Y49));
  sky130_fd_sc_hd__conb_1 conb_T24Y5 (.HI(tie_high_T24Y5), .LO(tie_low_T24Y5));
  sky130_fd_sc_hd__conb_1 conb_T24Y50 (.HI(tie_high_T24Y50), .LO(tie_low_T24Y50));
  sky130_fd_sc_hd__conb_1 conb_T24Y51 (.HI(tie_high_T24Y51), .LO(tie_low_T24Y51));
  sky130_fd_sc_hd__conb_1 conb_T24Y52 (.HI(tie_high_T24Y52), .LO(tie_low_T24Y52));
  sky130_fd_sc_hd__conb_1 conb_T24Y53 (.HI(tie_high_T24Y53), .LO(tie_low_T24Y53));
  sky130_fd_sc_hd__conb_1 conb_T24Y54 (.HI(tie_high_T24Y54), .LO(tie_low_T24Y54));
  sky130_fd_sc_hd__conb_1 conb_T24Y55 (.HI(tie_high_T24Y55), .LO(tie_low_T24Y55));
  sky130_fd_sc_hd__conb_1 conb_T24Y56 (.HI(tie_high_T24Y56), .LO(tie_low_T24Y56));
  sky130_fd_sc_hd__conb_1 conb_T24Y57 (.HI(tie_high_T24Y57), .LO(tie_low_T24Y57));
  sky130_fd_sc_hd__conb_1 conb_T24Y58 (.HI(tie_high_T24Y58), .LO(tie_low_T24Y58));
  sky130_fd_sc_hd__conb_1 conb_T24Y59 (.HI(tie_high_T24Y59), .LO(tie_low_T24Y59));
  sky130_fd_sc_hd__conb_1 conb_T24Y6 (.HI(tie_high_T24Y6), .LO(tie_low_T24Y6));
  sky130_fd_sc_hd__conb_1 conb_T24Y60 (.HI(tie_high_T24Y60), .LO(tie_low_T24Y60));
  sky130_fd_sc_hd__conb_1 conb_T24Y61 (.HI(tie_high_T24Y61), .LO(tie_low_T24Y61));
  sky130_fd_sc_hd__conb_1 conb_T24Y62 (.HI(tie_high_T24Y62), .LO(tie_low_T24Y62));
  sky130_fd_sc_hd__conb_1 conb_T24Y63 (.HI(tie_high_T24Y63), .LO(tie_low_T24Y63));
  sky130_fd_sc_hd__conb_1 conb_T24Y64 (.HI(tie_high_T24Y64), .LO(tie_low_T24Y64));
  sky130_fd_sc_hd__conb_1 conb_T24Y65 (.HI(tie_high_T24Y65), .LO(tie_low_T24Y65));
  sky130_fd_sc_hd__conb_1 conb_T24Y66 (.HI(tie_high_T24Y66), .LO(tie_low_T24Y66));
  sky130_fd_sc_hd__conb_1 conb_T24Y67 (.HI(tie_high_T24Y67), .LO(tie_low_T24Y67));
  sky130_fd_sc_hd__conb_1 conb_T24Y68 (.HI(tie_high_T24Y68), .LO(tie_low_T24Y68));
  sky130_fd_sc_hd__conb_1 conb_T24Y69 (.HI(tie_high_T24Y69), .LO(tie_low_T24Y69));
  sky130_fd_sc_hd__conb_1 conb_T24Y7 (.HI(tie_high_T24Y7), .LO(tie_low_T24Y7));
  sky130_fd_sc_hd__conb_1 conb_T24Y70 (.HI(tie_high_T24Y70), .LO(tie_low_T24Y70));
  sky130_fd_sc_hd__conb_1 conb_T24Y71 (.HI(tie_high_T24Y71), .LO(tie_low_T24Y71));
  sky130_fd_sc_hd__conb_1 conb_T24Y72 (.HI(tie_high_T24Y72), .LO(tie_low_T24Y72));
  sky130_fd_sc_hd__conb_1 conb_T24Y73 (.HI(tie_high_T24Y73), .LO(tie_low_T24Y73));
  sky130_fd_sc_hd__conb_1 conb_T24Y74 (.HI(tie_high_T24Y74), .LO(tie_low_T24Y74));
  sky130_fd_sc_hd__conb_1 conb_T24Y75 (.HI(tie_high_T24Y75), .LO(tie_low_T24Y75));
  sky130_fd_sc_hd__conb_1 conb_T24Y76 (.HI(tie_high_T24Y76), .LO(tie_low_T24Y76));
  sky130_fd_sc_hd__conb_1 conb_T24Y77 (.HI(tie_high_T24Y77), .LO(tie_low_T24Y77));
  sky130_fd_sc_hd__conb_1 conb_T24Y78 (.HI(tie_high_T24Y78), .LO(tie_low_T24Y78));
  sky130_fd_sc_hd__conb_1 conb_T24Y79 (.HI(tie_high_T24Y79), .LO(tie_low_T24Y79));
  sky130_fd_sc_hd__conb_1 conb_T24Y8 (.HI(tie_high_T24Y8), .LO(tie_low_T24Y8));
  sky130_fd_sc_hd__conb_1 conb_T24Y80 (.HI(tie_high_T24Y80), .LO(tie_low_T24Y80));
  sky130_fd_sc_hd__conb_1 conb_T24Y81 (.HI(tie_high_T24Y81), .LO(tie_low_T24Y81));
  sky130_fd_sc_hd__conb_1 conb_T24Y82 (.HI(tie_high_T24Y82), .LO(tie_low_T24Y82));
  sky130_fd_sc_hd__conb_1 conb_T24Y83 (.HI(tie_high_T24Y83), .LO(tie_low_T24Y83));
  sky130_fd_sc_hd__conb_1 conb_T24Y84 (.HI(tie_high_T24Y84), .LO(tie_low_T24Y84));
  sky130_fd_sc_hd__conb_1 conb_T24Y85 (.HI(tie_high_T24Y85), .LO(tie_low_T24Y85));
  sky130_fd_sc_hd__conb_1 conb_T24Y86 (.HI(tie_high_T24Y86), .LO(tie_low_T24Y86));
  sky130_fd_sc_hd__conb_1 conb_T24Y87 (.HI(tie_high_T24Y87), .LO(tie_low_T24Y87));
  sky130_fd_sc_hd__conb_1 conb_T24Y88 (.HI(tie_high_T24Y88), .LO(tie_low_T24Y88));
  sky130_fd_sc_hd__conb_1 conb_T24Y89 (.HI(tie_high_T24Y89), .LO(tie_low_T24Y89));
  sky130_fd_sc_hd__conb_1 conb_T24Y9 (.HI(tie_high_T24Y9), .LO(tie_low_T24Y9));
  sky130_fd_sc_hd__conb_1 conb_T25Y0 (.HI(tie_high_T25Y0), .LO(tie_low_T25Y0));
  sky130_fd_sc_hd__conb_1 conb_T25Y1 (.HI(tie_high_T25Y1), .LO(tie_low_T25Y1));
  sky130_fd_sc_hd__conb_1 conb_T25Y10 (.HI(tie_high_T25Y10), .LO(tie_low_T25Y10));
  sky130_fd_sc_hd__conb_1 conb_T25Y11 (.HI(tie_high_T25Y11), .LO(tie_low_T25Y11));
  sky130_fd_sc_hd__conb_1 conb_T25Y12 (.HI(tie_high_T25Y12), .LO(tie_low_T25Y12));
  sky130_fd_sc_hd__conb_1 conb_T25Y13 (.HI(tie_high_T25Y13), .LO(tie_low_T25Y13));
  sky130_fd_sc_hd__conb_1 conb_T25Y14 (.HI(tie_high_T25Y14), .LO(tie_low_T25Y14));
  sky130_fd_sc_hd__conb_1 conb_T25Y15 (.HI(tie_high_T25Y15), .LO(tie_low_T25Y15));
  sky130_fd_sc_hd__conb_1 conb_T25Y16 (.HI(tie_high_T25Y16), .LO(tie_low_T25Y16));
  sky130_fd_sc_hd__conb_1 conb_T25Y17 (.HI(tie_high_T25Y17), .LO(tie_low_T25Y17));
  sky130_fd_sc_hd__conb_1 conb_T25Y18 (.HI(tie_high_T25Y18), .LO(tie_low_T25Y18));
  sky130_fd_sc_hd__conb_1 conb_T25Y19 (.HI(tie_high_T25Y19), .LO(tie_low_T25Y19));
  sky130_fd_sc_hd__conb_1 conb_T25Y2 (.HI(tie_high_T25Y2), .LO(tie_low_T25Y2));
  sky130_fd_sc_hd__conb_1 conb_T25Y20 (.HI(tie_high_T25Y20), .LO(tie_low_T25Y20));
  sky130_fd_sc_hd__conb_1 conb_T25Y21 (.HI(tie_high_T25Y21), .LO(tie_low_T25Y21));
  sky130_fd_sc_hd__conb_1 conb_T25Y22 (.HI(tie_high_T25Y22), .LO(tie_low_T25Y22));
  sky130_fd_sc_hd__conb_1 conb_T25Y23 (.HI(tie_high_T25Y23), .LO(tie_low_T25Y23));
  sky130_fd_sc_hd__conb_1 conb_T25Y24 (.HI(tie_high_T25Y24), .LO(tie_low_T25Y24));
  sky130_fd_sc_hd__conb_1 conb_T25Y25 (.HI(tie_high_T25Y25), .LO(tie_low_T25Y25));
  sky130_fd_sc_hd__conb_1 conb_T25Y26 (.HI(tie_high_T25Y26), .LO(tie_low_T25Y26));
  sky130_fd_sc_hd__conb_1 conb_T25Y27 (.HI(tie_high_T25Y27), .LO(tie_low_T25Y27));
  sky130_fd_sc_hd__conb_1 conb_T25Y28 (.HI(tie_high_T25Y28), .LO(tie_low_T25Y28));
  sky130_fd_sc_hd__conb_1 conb_T25Y29 (.HI(tie_high_T25Y29), .LO(tie_low_T25Y29));
  sky130_fd_sc_hd__conb_1 conb_T25Y3 (.HI(tie_high_T25Y3), .LO(tie_low_T25Y3));
  sky130_fd_sc_hd__conb_1 conb_T25Y30 (.HI(tie_high_T25Y30), .LO(tie_low_T25Y30));
  sky130_fd_sc_hd__conb_1 conb_T25Y31 (.HI(tie_high_T25Y31), .LO(tie_low_T25Y31));
  sky130_fd_sc_hd__conb_1 conb_T25Y32 (.HI(tie_high_T25Y32), .LO(tie_low_T25Y32));
  sky130_fd_sc_hd__conb_1 conb_T25Y33 (.HI(tie_high_T25Y33), .LO(tie_low_T25Y33));
  sky130_fd_sc_hd__conb_1 conb_T25Y34 (.HI(tie_high_T25Y34), .LO(tie_low_T25Y34));
  sky130_fd_sc_hd__conb_1 conb_T25Y35 (.HI(tie_high_T25Y35), .LO(tie_low_T25Y35));
  sky130_fd_sc_hd__conb_1 conb_T25Y36 (.HI(tie_high_T25Y36), .LO(tie_low_T25Y36));
  sky130_fd_sc_hd__conb_1 conb_T25Y37 (.HI(tie_high_T25Y37), .LO(tie_low_T25Y37));
  sky130_fd_sc_hd__conb_1 conb_T25Y38 (.HI(tie_high_T25Y38), .LO(tie_low_T25Y38));
  sky130_fd_sc_hd__conb_1 conb_T25Y39 (.HI(tie_high_T25Y39), .LO(tie_low_T25Y39));
  sky130_fd_sc_hd__conb_1 conb_T25Y4 (.HI(tie_high_T25Y4), .LO(tie_low_T25Y4));
  sky130_fd_sc_hd__conb_1 conb_T25Y40 (.HI(tie_high_T25Y40), .LO(tie_low_T25Y40));
  sky130_fd_sc_hd__conb_1 conb_T25Y41 (.HI(tie_high_T25Y41), .LO(tie_low_T25Y41));
  sky130_fd_sc_hd__conb_1 conb_T25Y42 (.HI(tie_high_T25Y42), .LO(tie_low_T25Y42));
  sky130_fd_sc_hd__conb_1 conb_T25Y43 (.HI(tie_high_T25Y43), .LO(tie_low_T25Y43));
  sky130_fd_sc_hd__conb_1 conb_T25Y44 (.HI(tie_high_T25Y44), .LO(tie_low_T25Y44));
  sky130_fd_sc_hd__conb_1 conb_T25Y45 (.HI(tie_high_T25Y45), .LO(tie_low_T25Y45));
  sky130_fd_sc_hd__conb_1 conb_T25Y46 (.HI(tie_high_T25Y46), .LO(tie_low_T25Y46));
  sky130_fd_sc_hd__conb_1 conb_T25Y47 (.HI(tie_high_T25Y47), .LO(tie_low_T25Y47));
  sky130_fd_sc_hd__conb_1 conb_T25Y48 (.HI(tie_high_T25Y48), .LO(tie_low_T25Y48));
  sky130_fd_sc_hd__conb_1 conb_T25Y49 (.HI(tie_high_T25Y49), .LO(tie_low_T25Y49));
  sky130_fd_sc_hd__conb_1 conb_T25Y5 (.HI(tie_high_T25Y5), .LO(tie_low_T25Y5));
  sky130_fd_sc_hd__conb_1 conb_T25Y50 (.HI(tie_high_T25Y50), .LO(tie_low_T25Y50));
  sky130_fd_sc_hd__conb_1 conb_T25Y51 (.HI(tie_high_T25Y51), .LO(tie_low_T25Y51));
  sky130_fd_sc_hd__conb_1 conb_T25Y52 (.HI(tie_high_T25Y52), .LO(tie_low_T25Y52));
  sky130_fd_sc_hd__conb_1 conb_T25Y53 (.HI(tie_high_T25Y53), .LO(tie_low_T25Y53));
  sky130_fd_sc_hd__conb_1 conb_T25Y54 (.HI(tie_high_T25Y54), .LO(tie_low_T25Y54));
  sky130_fd_sc_hd__conb_1 conb_T25Y55 (.HI(tie_high_T25Y55), .LO(tie_low_T25Y55));
  sky130_fd_sc_hd__conb_1 conb_T25Y56 (.HI(tie_high_T25Y56), .LO(tie_low_T25Y56));
  sky130_fd_sc_hd__conb_1 conb_T25Y57 (.HI(tie_high_T25Y57), .LO(tie_low_T25Y57));
  sky130_fd_sc_hd__conb_1 conb_T25Y58 (.HI(tie_high_T25Y58), .LO(tie_low_T25Y58));
  sky130_fd_sc_hd__conb_1 conb_T25Y59 (.HI(tie_high_T25Y59), .LO(tie_low_T25Y59));
  sky130_fd_sc_hd__conb_1 conb_T25Y6 (.HI(tie_high_T25Y6), .LO(tie_low_T25Y6));
  sky130_fd_sc_hd__conb_1 conb_T25Y60 (.HI(tie_high_T25Y60), .LO(tie_low_T25Y60));
  sky130_fd_sc_hd__conb_1 conb_T25Y61 (.HI(tie_high_T25Y61), .LO(tie_low_T25Y61));
  sky130_fd_sc_hd__conb_1 conb_T25Y62 (.HI(tie_high_T25Y62), .LO(tie_low_T25Y62));
  sky130_fd_sc_hd__conb_1 conb_T25Y63 (.HI(tie_high_T25Y63), .LO(tie_low_T25Y63));
  sky130_fd_sc_hd__conb_1 conb_T25Y64 (.HI(tie_high_T25Y64), .LO(tie_low_T25Y64));
  sky130_fd_sc_hd__conb_1 conb_T25Y65 (.HI(tie_high_T25Y65), .LO(tie_low_T25Y65));
  sky130_fd_sc_hd__conb_1 conb_T25Y66 (.HI(tie_high_T25Y66), .LO(tie_low_T25Y66));
  sky130_fd_sc_hd__conb_1 conb_T25Y67 (.HI(tie_high_T25Y67), .LO(tie_low_T25Y67));
  sky130_fd_sc_hd__conb_1 conb_T25Y68 (.HI(tie_high_T25Y68), .LO(tie_low_T25Y68));
  sky130_fd_sc_hd__conb_1 conb_T25Y69 (.HI(tie_high_T25Y69), .LO(tie_low_T25Y69));
  sky130_fd_sc_hd__conb_1 conb_T25Y7 (.HI(tie_high_T25Y7), .LO(tie_low_T25Y7));
  sky130_fd_sc_hd__conb_1 conb_T25Y70 (.HI(tie_high_T25Y70), .LO(tie_low_T25Y70));
  sky130_fd_sc_hd__conb_1 conb_T25Y71 (.HI(tie_high_T25Y71), .LO(tie_low_T25Y71));
  sky130_fd_sc_hd__conb_1 conb_T25Y72 (.HI(tie_high_T25Y72), .LO(tie_low_T25Y72));
  sky130_fd_sc_hd__conb_1 conb_T25Y73 (.HI(tie_high_T25Y73), .LO(tie_low_T25Y73));
  sky130_fd_sc_hd__conb_1 conb_T25Y74 (.HI(tie_high_T25Y74), .LO(tie_low_T25Y74));
  sky130_fd_sc_hd__conb_1 conb_T25Y75 (.HI(tie_high_T25Y75), .LO(tie_low_T25Y75));
  sky130_fd_sc_hd__conb_1 conb_T25Y76 (.HI(tie_high_T25Y76), .LO(tie_low_T25Y76));
  sky130_fd_sc_hd__conb_1 conb_T25Y77 (.HI(tie_high_T25Y77), .LO(tie_low_T25Y77));
  sky130_fd_sc_hd__conb_1 conb_T25Y78 (.HI(tie_high_T25Y78), .LO(tie_low_T25Y78));
  sky130_fd_sc_hd__conb_1 conb_T25Y79 (.HI(tie_high_T25Y79), .LO(tie_low_T25Y79));
  sky130_fd_sc_hd__conb_1 conb_T25Y8 (.HI(tie_high_T25Y8), .LO(tie_low_T25Y8));
  sky130_fd_sc_hd__conb_1 conb_T25Y80 (.HI(tie_high_T25Y80), .LO(tie_low_T25Y80));
  sky130_fd_sc_hd__conb_1 conb_T25Y81 (.HI(tie_high_T25Y81), .LO(tie_low_T25Y81));
  sky130_fd_sc_hd__conb_1 conb_T25Y82 (.HI(tie_high_T25Y82), .LO(tie_low_T25Y82));
  sky130_fd_sc_hd__conb_1 conb_T25Y83 (.HI(tie_high_T25Y83), .LO(tie_low_T25Y83));
  sky130_fd_sc_hd__conb_1 conb_T25Y84 (.HI(tie_high_T25Y84), .LO(tie_low_T25Y84));
  sky130_fd_sc_hd__conb_1 conb_T25Y85 (.HI(tie_high_T25Y85), .LO(tie_low_T25Y85));
  sky130_fd_sc_hd__conb_1 conb_T25Y86 (.HI(tie_high_T25Y86), .LO(tie_low_T25Y86));
  sky130_fd_sc_hd__conb_1 conb_T25Y87 (.HI(tie_high_T25Y87), .LO(tie_low_T25Y87));
  sky130_fd_sc_hd__conb_1 conb_T25Y88 (.HI(tie_high_T25Y88), .LO(tie_low_T25Y88));
  sky130_fd_sc_hd__conb_1 conb_T25Y89 (.HI(tie_high_T25Y89), .LO(tie_low_T25Y89));
  sky130_fd_sc_hd__conb_1 conb_T25Y9 (.HI(tie_high_T25Y9), .LO(tie_low_T25Y9));
  sky130_fd_sc_hd__conb_1 conb_T26Y0 (.HI(tie_high_T26Y0), .LO(tie_low_T26Y0));
  sky130_fd_sc_hd__conb_1 conb_T26Y1 (.HI(tie_high_T26Y1), .LO(tie_low_T26Y1));
  sky130_fd_sc_hd__conb_1 conb_T26Y10 (.HI(tie_high_T26Y10), .LO(tie_low_T26Y10));
  sky130_fd_sc_hd__conb_1 conb_T26Y11 (.HI(tie_high_T26Y11), .LO(tie_low_T26Y11));
  sky130_fd_sc_hd__conb_1 conb_T26Y12 (.HI(tie_high_T26Y12), .LO(tie_low_T26Y12));
  sky130_fd_sc_hd__conb_1 conb_T26Y13 (.HI(tie_high_T26Y13), .LO(tie_low_T26Y13));
  sky130_fd_sc_hd__conb_1 conb_T26Y14 (.HI(tie_high_T26Y14), .LO(tie_low_T26Y14));
  sky130_fd_sc_hd__conb_1 conb_T26Y15 (.HI(tie_high_T26Y15), .LO(tie_low_T26Y15));
  sky130_fd_sc_hd__conb_1 conb_T26Y16 (.HI(tie_high_T26Y16), .LO(tie_low_T26Y16));
  sky130_fd_sc_hd__conb_1 conb_T26Y17 (.HI(tie_high_T26Y17), .LO(tie_low_T26Y17));
  sky130_fd_sc_hd__conb_1 conb_T26Y18 (.HI(tie_high_T26Y18), .LO(tie_low_T26Y18));
  sky130_fd_sc_hd__conb_1 conb_T26Y19 (.HI(tie_high_T26Y19), .LO(tie_low_T26Y19));
  sky130_fd_sc_hd__conb_1 conb_T26Y2 (.HI(tie_high_T26Y2), .LO(tie_low_T26Y2));
  sky130_fd_sc_hd__conb_1 conb_T26Y20 (.HI(tie_high_T26Y20), .LO(tie_low_T26Y20));
  sky130_fd_sc_hd__conb_1 conb_T26Y21 (.HI(tie_high_T26Y21), .LO(tie_low_T26Y21));
  sky130_fd_sc_hd__conb_1 conb_T26Y22 (.HI(tie_high_T26Y22), .LO(tie_low_T26Y22));
  sky130_fd_sc_hd__conb_1 conb_T26Y23 (.HI(tie_high_T26Y23), .LO(tie_low_T26Y23));
  sky130_fd_sc_hd__conb_1 conb_T26Y24 (.HI(tie_high_T26Y24), .LO(tie_low_T26Y24));
  sky130_fd_sc_hd__conb_1 conb_T26Y25 (.HI(tie_high_T26Y25), .LO(tie_low_T26Y25));
  sky130_fd_sc_hd__conb_1 conb_T26Y26 (.HI(tie_high_T26Y26), .LO(tie_low_T26Y26));
  sky130_fd_sc_hd__conb_1 conb_T26Y27 (.HI(tie_high_T26Y27), .LO(tie_low_T26Y27));
  sky130_fd_sc_hd__conb_1 conb_T26Y28 (.HI(tie_high_T26Y28), .LO(tie_low_T26Y28));
  sky130_fd_sc_hd__conb_1 conb_T26Y29 (.HI(tie_high_T26Y29), .LO(tie_low_T26Y29));
  sky130_fd_sc_hd__conb_1 conb_T26Y3 (.HI(tie_high_T26Y3), .LO(tie_low_T26Y3));
  sky130_fd_sc_hd__conb_1 conb_T26Y30 (.HI(tie_high_T26Y30), .LO(tie_low_T26Y30));
  sky130_fd_sc_hd__conb_1 conb_T26Y31 (.HI(tie_high_T26Y31), .LO(tie_low_T26Y31));
  sky130_fd_sc_hd__conb_1 conb_T26Y32 (.HI(tie_high_T26Y32), .LO(tie_low_T26Y32));
  sky130_fd_sc_hd__conb_1 conb_T26Y33 (.HI(tie_high_T26Y33), .LO(tie_low_T26Y33));
  sky130_fd_sc_hd__conb_1 conb_T26Y34 (.HI(tie_high_T26Y34), .LO(tie_low_T26Y34));
  sky130_fd_sc_hd__conb_1 conb_T26Y35 (.HI(tie_high_T26Y35), .LO(tie_low_T26Y35));
  sky130_fd_sc_hd__conb_1 conb_T26Y36 (.HI(tie_high_T26Y36), .LO(tie_low_T26Y36));
  sky130_fd_sc_hd__conb_1 conb_T26Y37 (.HI(tie_high_T26Y37), .LO(tie_low_T26Y37));
  sky130_fd_sc_hd__conb_1 conb_T26Y38 (.HI(tie_high_T26Y38), .LO(tie_low_T26Y38));
  sky130_fd_sc_hd__conb_1 conb_T26Y39 (.HI(tie_high_T26Y39), .LO(tie_low_T26Y39));
  sky130_fd_sc_hd__conb_1 conb_T26Y4 (.HI(tie_high_T26Y4), .LO(tie_low_T26Y4));
  sky130_fd_sc_hd__conb_1 conb_T26Y40 (.HI(tie_high_T26Y40), .LO(tie_low_T26Y40));
  sky130_fd_sc_hd__conb_1 conb_T26Y41 (.HI(tie_high_T26Y41), .LO(tie_low_T26Y41));
  sky130_fd_sc_hd__conb_1 conb_T26Y42 (.HI(tie_high_T26Y42), .LO(tie_low_T26Y42));
  sky130_fd_sc_hd__conb_1 conb_T26Y43 (.HI(tie_high_T26Y43), .LO(tie_low_T26Y43));
  sky130_fd_sc_hd__conb_1 conb_T26Y44 (.HI(tie_high_T26Y44), .LO(tie_low_T26Y44));
  sky130_fd_sc_hd__conb_1 conb_T26Y45 (.HI(tie_high_T26Y45), .LO(tie_low_T26Y45));
  sky130_fd_sc_hd__conb_1 conb_T26Y46 (.HI(tie_high_T26Y46), .LO(tie_low_T26Y46));
  sky130_fd_sc_hd__conb_1 conb_T26Y47 (.HI(tie_high_T26Y47), .LO(tie_low_T26Y47));
  sky130_fd_sc_hd__conb_1 conb_T26Y48 (.HI(tie_high_T26Y48), .LO(tie_low_T26Y48));
  sky130_fd_sc_hd__conb_1 conb_T26Y49 (.HI(tie_high_T26Y49), .LO(tie_low_T26Y49));
  sky130_fd_sc_hd__conb_1 conb_T26Y5 (.HI(tie_high_T26Y5), .LO(tie_low_T26Y5));
  sky130_fd_sc_hd__conb_1 conb_T26Y50 (.HI(tie_high_T26Y50), .LO(tie_low_T26Y50));
  sky130_fd_sc_hd__conb_1 conb_T26Y51 (.HI(tie_high_T26Y51), .LO(tie_low_T26Y51));
  sky130_fd_sc_hd__conb_1 conb_T26Y52 (.HI(tie_high_T26Y52), .LO(tie_low_T26Y52));
  sky130_fd_sc_hd__conb_1 conb_T26Y53 (.HI(tie_high_T26Y53), .LO(tie_low_T26Y53));
  sky130_fd_sc_hd__conb_1 conb_T26Y54 (.HI(tie_high_T26Y54), .LO(tie_low_T26Y54));
  sky130_fd_sc_hd__conb_1 conb_T26Y55 (.HI(tie_high_T26Y55), .LO(tie_low_T26Y55));
  sky130_fd_sc_hd__conb_1 conb_T26Y56 (.HI(tie_high_T26Y56), .LO(tie_low_T26Y56));
  sky130_fd_sc_hd__conb_1 conb_T26Y57 (.HI(tie_high_T26Y57), .LO(tie_low_T26Y57));
  sky130_fd_sc_hd__conb_1 conb_T26Y58 (.HI(tie_high_T26Y58), .LO(tie_low_T26Y58));
  sky130_fd_sc_hd__conb_1 conb_T26Y59 (.HI(tie_high_T26Y59), .LO(tie_low_T26Y59));
  sky130_fd_sc_hd__conb_1 conb_T26Y6 (.HI(tie_high_T26Y6), .LO(tie_low_T26Y6));
  sky130_fd_sc_hd__conb_1 conb_T26Y60 (.HI(tie_high_T26Y60), .LO(tie_low_T26Y60));
  sky130_fd_sc_hd__conb_1 conb_T26Y61 (.HI(tie_high_T26Y61), .LO(tie_low_T26Y61));
  sky130_fd_sc_hd__conb_1 conb_T26Y62 (.HI(tie_high_T26Y62), .LO(tie_low_T26Y62));
  sky130_fd_sc_hd__conb_1 conb_T26Y63 (.HI(tie_high_T26Y63), .LO(tie_low_T26Y63));
  sky130_fd_sc_hd__conb_1 conb_T26Y64 (.HI(tie_high_T26Y64), .LO(tie_low_T26Y64));
  sky130_fd_sc_hd__conb_1 conb_T26Y65 (.HI(tie_high_T26Y65), .LO(tie_low_T26Y65));
  sky130_fd_sc_hd__conb_1 conb_T26Y66 (.HI(tie_high_T26Y66), .LO(tie_low_T26Y66));
  sky130_fd_sc_hd__conb_1 conb_T26Y67 (.HI(tie_high_T26Y67), .LO(tie_low_T26Y67));
  sky130_fd_sc_hd__conb_1 conb_T26Y68 (.HI(tie_high_T26Y68), .LO(tie_low_T26Y68));
  sky130_fd_sc_hd__conb_1 conb_T26Y69 (.HI(tie_high_T26Y69), .LO(tie_low_T26Y69));
  sky130_fd_sc_hd__conb_1 conb_T26Y7 (.HI(tie_high_T26Y7), .LO(tie_low_T26Y7));
  sky130_fd_sc_hd__conb_1 conb_T26Y70 (.HI(tie_high_T26Y70), .LO(tie_low_T26Y70));
  sky130_fd_sc_hd__conb_1 conb_T26Y71 (.HI(tie_high_T26Y71), .LO(tie_low_T26Y71));
  sky130_fd_sc_hd__conb_1 conb_T26Y72 (.HI(tie_high_T26Y72), .LO(tie_low_T26Y72));
  sky130_fd_sc_hd__conb_1 conb_T26Y73 (.HI(tie_high_T26Y73), .LO(tie_low_T26Y73));
  sky130_fd_sc_hd__conb_1 conb_T26Y74 (.HI(tie_high_T26Y74), .LO(tie_low_T26Y74));
  sky130_fd_sc_hd__conb_1 conb_T26Y75 (.HI(tie_high_T26Y75), .LO(tie_low_T26Y75));
  sky130_fd_sc_hd__conb_1 conb_T26Y76 (.HI(tie_high_T26Y76), .LO(tie_low_T26Y76));
  sky130_fd_sc_hd__conb_1 conb_T26Y77 (.HI(tie_high_T26Y77), .LO(tie_low_T26Y77));
  sky130_fd_sc_hd__conb_1 conb_T26Y78 (.HI(tie_high_T26Y78), .LO(tie_low_T26Y78));
  sky130_fd_sc_hd__conb_1 conb_T26Y79 (.HI(tie_high_T26Y79), .LO(tie_low_T26Y79));
  sky130_fd_sc_hd__conb_1 conb_T26Y8 (.HI(tie_high_T26Y8), .LO(tie_low_T26Y8));
  sky130_fd_sc_hd__conb_1 conb_T26Y80 (.HI(tie_high_T26Y80), .LO(tie_low_T26Y80));
  sky130_fd_sc_hd__conb_1 conb_T26Y81 (.HI(tie_high_T26Y81), .LO(tie_low_T26Y81));
  sky130_fd_sc_hd__conb_1 conb_T26Y82 (.HI(tie_high_T26Y82), .LO(tie_low_T26Y82));
  sky130_fd_sc_hd__conb_1 conb_T26Y83 (.HI(tie_high_T26Y83), .LO(tie_low_T26Y83));
  sky130_fd_sc_hd__conb_1 conb_T26Y84 (.HI(tie_high_T26Y84), .LO(tie_low_T26Y84));
  sky130_fd_sc_hd__conb_1 conb_T26Y85 (.HI(tie_high_T26Y85), .LO(tie_low_T26Y85));
  sky130_fd_sc_hd__conb_1 conb_T26Y86 (.HI(tie_high_T26Y86), .LO(tie_low_T26Y86));
  sky130_fd_sc_hd__conb_1 conb_T26Y87 (.HI(tie_high_T26Y87), .LO(tie_low_T26Y87));
  sky130_fd_sc_hd__conb_1 conb_T26Y88 (.HI(tie_high_T26Y88), .LO(tie_low_T26Y88));
  sky130_fd_sc_hd__conb_1 conb_T26Y89 (.HI(tie_high_T26Y89), .LO(tie_low_T26Y89));
  sky130_fd_sc_hd__conb_1 conb_T26Y9 (.HI(tie_high_T26Y9), .LO(tie_low_T26Y9));
  sky130_fd_sc_hd__conb_1 conb_T27Y0 (.HI(tie_high_T27Y0), .LO(tie_low_T27Y0));
  sky130_fd_sc_hd__conb_1 conb_T27Y1 (.HI(tie_high_T27Y1), .LO(tie_low_T27Y1));
  sky130_fd_sc_hd__conb_1 conb_T27Y10 (.HI(tie_high_T27Y10), .LO(tie_low_T27Y10));
  sky130_fd_sc_hd__conb_1 conb_T27Y11 (.HI(tie_high_T27Y11), .LO(tie_low_T27Y11));
  sky130_fd_sc_hd__conb_1 conb_T27Y12 (.HI(tie_high_T27Y12), .LO(tie_low_T27Y12));
  sky130_fd_sc_hd__conb_1 conb_T27Y13 (.HI(tie_high_T27Y13), .LO(tie_low_T27Y13));
  sky130_fd_sc_hd__conb_1 conb_T27Y14 (.HI(tie_high_T27Y14), .LO(tie_low_T27Y14));
  sky130_fd_sc_hd__conb_1 conb_T27Y15 (.HI(tie_high_T27Y15), .LO(tie_low_T27Y15));
  sky130_fd_sc_hd__conb_1 conb_T27Y16 (.HI(tie_high_T27Y16), .LO(tie_low_T27Y16));
  sky130_fd_sc_hd__conb_1 conb_T27Y17 (.HI(tie_high_T27Y17), .LO(tie_low_T27Y17));
  sky130_fd_sc_hd__conb_1 conb_T27Y18 (.HI(tie_high_T27Y18), .LO(tie_low_T27Y18));
  sky130_fd_sc_hd__conb_1 conb_T27Y19 (.HI(tie_high_T27Y19), .LO(tie_low_T27Y19));
  sky130_fd_sc_hd__conb_1 conb_T27Y2 (.HI(tie_high_T27Y2), .LO(tie_low_T27Y2));
  sky130_fd_sc_hd__conb_1 conb_T27Y20 (.HI(tie_high_T27Y20), .LO(tie_low_T27Y20));
  sky130_fd_sc_hd__conb_1 conb_T27Y21 (.HI(tie_high_T27Y21), .LO(tie_low_T27Y21));
  sky130_fd_sc_hd__conb_1 conb_T27Y22 (.HI(tie_high_T27Y22), .LO(tie_low_T27Y22));
  sky130_fd_sc_hd__conb_1 conb_T27Y23 (.HI(tie_high_T27Y23), .LO(tie_low_T27Y23));
  sky130_fd_sc_hd__conb_1 conb_T27Y24 (.HI(tie_high_T27Y24), .LO(tie_low_T27Y24));
  sky130_fd_sc_hd__conb_1 conb_T27Y25 (.HI(tie_high_T27Y25), .LO(tie_low_T27Y25));
  sky130_fd_sc_hd__conb_1 conb_T27Y26 (.HI(tie_high_T27Y26), .LO(tie_low_T27Y26));
  sky130_fd_sc_hd__conb_1 conb_T27Y27 (.HI(tie_high_T27Y27), .LO(tie_low_T27Y27));
  sky130_fd_sc_hd__conb_1 conb_T27Y28 (.HI(tie_high_T27Y28), .LO(tie_low_T27Y28));
  sky130_fd_sc_hd__conb_1 conb_T27Y29 (.HI(tie_high_T27Y29), .LO(tie_low_T27Y29));
  sky130_fd_sc_hd__conb_1 conb_T27Y3 (.HI(tie_high_T27Y3), .LO(tie_low_T27Y3));
  sky130_fd_sc_hd__conb_1 conb_T27Y30 (.HI(tie_high_T27Y30), .LO(tie_low_T27Y30));
  sky130_fd_sc_hd__conb_1 conb_T27Y31 (.HI(tie_high_T27Y31), .LO(tie_low_T27Y31));
  sky130_fd_sc_hd__conb_1 conb_T27Y32 (.HI(tie_high_T27Y32), .LO(tie_low_T27Y32));
  sky130_fd_sc_hd__conb_1 conb_T27Y33 (.HI(tie_high_T27Y33), .LO(tie_low_T27Y33));
  sky130_fd_sc_hd__conb_1 conb_T27Y34 (.HI(tie_high_T27Y34), .LO(tie_low_T27Y34));
  sky130_fd_sc_hd__conb_1 conb_T27Y35 (.HI(tie_high_T27Y35), .LO(tie_low_T27Y35));
  sky130_fd_sc_hd__conb_1 conb_T27Y36 (.HI(tie_high_T27Y36), .LO(tie_low_T27Y36));
  sky130_fd_sc_hd__conb_1 conb_T27Y37 (.HI(tie_high_T27Y37), .LO(tie_low_T27Y37));
  sky130_fd_sc_hd__conb_1 conb_T27Y38 (.HI(tie_high_T27Y38), .LO(tie_low_T27Y38));
  sky130_fd_sc_hd__conb_1 conb_T27Y39 (.HI(tie_high_T27Y39), .LO(tie_low_T27Y39));
  sky130_fd_sc_hd__conb_1 conb_T27Y4 (.HI(tie_high_T27Y4), .LO(tie_low_T27Y4));
  sky130_fd_sc_hd__conb_1 conb_T27Y40 (.HI(tie_high_T27Y40), .LO(tie_low_T27Y40));
  sky130_fd_sc_hd__conb_1 conb_T27Y41 (.HI(tie_high_T27Y41), .LO(tie_low_T27Y41));
  sky130_fd_sc_hd__conb_1 conb_T27Y42 (.HI(tie_high_T27Y42), .LO(tie_low_T27Y42));
  sky130_fd_sc_hd__conb_1 conb_T27Y43 (.HI(tie_high_T27Y43), .LO(tie_low_T27Y43));
  sky130_fd_sc_hd__conb_1 conb_T27Y44 (.HI(tie_high_T27Y44), .LO(tie_low_T27Y44));
  sky130_fd_sc_hd__conb_1 conb_T27Y45 (.HI(tie_high_T27Y45), .LO(tie_low_T27Y45));
  sky130_fd_sc_hd__conb_1 conb_T27Y46 (.HI(tie_high_T27Y46), .LO(tie_low_T27Y46));
  sky130_fd_sc_hd__conb_1 conb_T27Y47 (.HI(tie_high_T27Y47), .LO(tie_low_T27Y47));
  sky130_fd_sc_hd__conb_1 conb_T27Y48 (.HI(tie_high_T27Y48), .LO(tie_low_T27Y48));
  sky130_fd_sc_hd__conb_1 conb_T27Y49 (.HI(tie_high_T27Y49), .LO(tie_low_T27Y49));
  sky130_fd_sc_hd__conb_1 conb_T27Y5 (.HI(tie_high_T27Y5), .LO(tie_low_T27Y5));
  sky130_fd_sc_hd__conb_1 conb_T27Y50 (.HI(tie_high_T27Y50), .LO(tie_low_T27Y50));
  sky130_fd_sc_hd__conb_1 conb_T27Y51 (.HI(tie_high_T27Y51), .LO(tie_low_T27Y51));
  sky130_fd_sc_hd__conb_1 conb_T27Y52 (.HI(tie_high_T27Y52), .LO(tie_low_T27Y52));
  sky130_fd_sc_hd__conb_1 conb_T27Y53 (.HI(tie_high_T27Y53), .LO(tie_low_T27Y53));
  sky130_fd_sc_hd__conb_1 conb_T27Y54 (.HI(tie_high_T27Y54), .LO(tie_low_T27Y54));
  sky130_fd_sc_hd__conb_1 conb_T27Y55 (.HI(tie_high_T27Y55), .LO(tie_low_T27Y55));
  sky130_fd_sc_hd__conb_1 conb_T27Y56 (.HI(tie_high_T27Y56), .LO(tie_low_T27Y56));
  sky130_fd_sc_hd__conb_1 conb_T27Y57 (.HI(tie_high_T27Y57), .LO(tie_low_T27Y57));
  sky130_fd_sc_hd__conb_1 conb_T27Y58 (.HI(tie_high_T27Y58), .LO(tie_low_T27Y58));
  sky130_fd_sc_hd__conb_1 conb_T27Y59 (.HI(tie_high_T27Y59), .LO(tie_low_T27Y59));
  sky130_fd_sc_hd__conb_1 conb_T27Y6 (.HI(tie_high_T27Y6), .LO(tie_low_T27Y6));
  sky130_fd_sc_hd__conb_1 conb_T27Y60 (.HI(tie_high_T27Y60), .LO(tie_low_T27Y60));
  sky130_fd_sc_hd__conb_1 conb_T27Y61 (.HI(tie_high_T27Y61), .LO(tie_low_T27Y61));
  sky130_fd_sc_hd__conb_1 conb_T27Y62 (.HI(tie_high_T27Y62), .LO(tie_low_T27Y62));
  sky130_fd_sc_hd__conb_1 conb_T27Y63 (.HI(tie_high_T27Y63), .LO(tie_low_T27Y63));
  sky130_fd_sc_hd__conb_1 conb_T27Y64 (.HI(tie_high_T27Y64), .LO(tie_low_T27Y64));
  sky130_fd_sc_hd__conb_1 conb_T27Y65 (.HI(tie_high_T27Y65), .LO(tie_low_T27Y65));
  sky130_fd_sc_hd__conb_1 conb_T27Y66 (.HI(tie_high_T27Y66), .LO(tie_low_T27Y66));
  sky130_fd_sc_hd__conb_1 conb_T27Y67 (.HI(tie_high_T27Y67), .LO(tie_low_T27Y67));
  sky130_fd_sc_hd__conb_1 conb_T27Y68 (.HI(tie_high_T27Y68), .LO(tie_low_T27Y68));
  sky130_fd_sc_hd__conb_1 conb_T27Y69 (.HI(tie_high_T27Y69), .LO(tie_low_T27Y69));
  sky130_fd_sc_hd__conb_1 conb_T27Y7 (.HI(tie_high_T27Y7), .LO(tie_low_T27Y7));
  sky130_fd_sc_hd__conb_1 conb_T27Y70 (.HI(tie_high_T27Y70), .LO(tie_low_T27Y70));
  sky130_fd_sc_hd__conb_1 conb_T27Y71 (.HI(tie_high_T27Y71), .LO(tie_low_T27Y71));
  sky130_fd_sc_hd__conb_1 conb_T27Y72 (.HI(tie_high_T27Y72), .LO(tie_low_T27Y72));
  sky130_fd_sc_hd__conb_1 conb_T27Y73 (.HI(tie_high_T27Y73), .LO(tie_low_T27Y73));
  sky130_fd_sc_hd__conb_1 conb_T27Y74 (.HI(tie_high_T27Y74), .LO(tie_low_T27Y74));
  sky130_fd_sc_hd__conb_1 conb_T27Y75 (.HI(tie_high_T27Y75), .LO(tie_low_T27Y75));
  sky130_fd_sc_hd__conb_1 conb_T27Y76 (.HI(tie_high_T27Y76), .LO(tie_low_T27Y76));
  sky130_fd_sc_hd__conb_1 conb_T27Y77 (.HI(tie_high_T27Y77), .LO(tie_low_T27Y77));
  sky130_fd_sc_hd__conb_1 conb_T27Y78 (.HI(tie_high_T27Y78), .LO(tie_low_T27Y78));
  sky130_fd_sc_hd__conb_1 conb_T27Y79 (.HI(tie_high_T27Y79), .LO(tie_low_T27Y79));
  sky130_fd_sc_hd__conb_1 conb_T27Y8 (.HI(tie_high_T27Y8), .LO(tie_low_T27Y8));
  sky130_fd_sc_hd__conb_1 conb_T27Y80 (.HI(tie_high_T27Y80), .LO(tie_low_T27Y80));
  sky130_fd_sc_hd__conb_1 conb_T27Y81 (.HI(tie_high_T27Y81), .LO(tie_low_T27Y81));
  sky130_fd_sc_hd__conb_1 conb_T27Y82 (.HI(tie_high_T27Y82), .LO(tie_low_T27Y82));
  sky130_fd_sc_hd__conb_1 conb_T27Y83 (.HI(tie_high_T27Y83), .LO(tie_low_T27Y83));
  sky130_fd_sc_hd__conb_1 conb_T27Y84 (.HI(tie_high_T27Y84), .LO(tie_low_T27Y84));
  sky130_fd_sc_hd__conb_1 conb_T27Y85 (.HI(tie_high_T27Y85), .LO(tie_low_T27Y85));
  sky130_fd_sc_hd__conb_1 conb_T27Y86 (.HI(tie_high_T27Y86), .LO(tie_low_T27Y86));
  sky130_fd_sc_hd__conb_1 conb_T27Y87 (.HI(tie_high_T27Y87), .LO(tie_low_T27Y87));
  sky130_fd_sc_hd__conb_1 conb_T27Y88 (.HI(tie_high_T27Y88), .LO(tie_low_T27Y88));
  sky130_fd_sc_hd__conb_1 conb_T27Y89 (.HI(tie_high_T27Y89), .LO(tie_low_T27Y89));
  sky130_fd_sc_hd__conb_1 conb_T27Y9 (.HI(tie_high_T27Y9), .LO(tie_low_T27Y9));
  sky130_fd_sc_hd__conb_1 conb_T28Y0 (.HI(tie_high_T28Y0), .LO(tie_low_T28Y0));
  sky130_fd_sc_hd__conb_1 conb_T28Y1 (.HI(tie_high_T28Y1), .LO(tie_low_T28Y1));
  sky130_fd_sc_hd__conb_1 conb_T28Y10 (.HI(tie_high_T28Y10), .LO(tie_low_T28Y10));
  sky130_fd_sc_hd__conb_1 conb_T28Y11 (.HI(tie_high_T28Y11), .LO(tie_low_T28Y11));
  sky130_fd_sc_hd__conb_1 conb_T28Y12 (.HI(tie_high_T28Y12), .LO(tie_low_T28Y12));
  sky130_fd_sc_hd__conb_1 conb_T28Y13 (.HI(tie_high_T28Y13), .LO(tie_low_T28Y13));
  sky130_fd_sc_hd__conb_1 conb_T28Y14 (.HI(tie_high_T28Y14), .LO(tie_low_T28Y14));
  sky130_fd_sc_hd__conb_1 conb_T28Y15 (.HI(tie_high_T28Y15), .LO(tie_low_T28Y15));
  sky130_fd_sc_hd__conb_1 conb_T28Y16 (.HI(tie_high_T28Y16), .LO(tie_low_T28Y16));
  sky130_fd_sc_hd__conb_1 conb_T28Y17 (.HI(tie_high_T28Y17), .LO(tie_low_T28Y17));
  sky130_fd_sc_hd__conb_1 conb_T28Y18 (.HI(tie_high_T28Y18), .LO(tie_low_T28Y18));
  sky130_fd_sc_hd__conb_1 conb_T28Y19 (.HI(tie_high_T28Y19), .LO(tie_low_T28Y19));
  sky130_fd_sc_hd__conb_1 conb_T28Y2 (.HI(tie_high_T28Y2), .LO(tie_low_T28Y2));
  sky130_fd_sc_hd__conb_1 conb_T28Y20 (.HI(tie_high_T28Y20), .LO(tie_low_T28Y20));
  sky130_fd_sc_hd__conb_1 conb_T28Y21 (.HI(tie_high_T28Y21), .LO(tie_low_T28Y21));
  sky130_fd_sc_hd__conb_1 conb_T28Y22 (.HI(tie_high_T28Y22), .LO(tie_low_T28Y22));
  sky130_fd_sc_hd__conb_1 conb_T28Y23 (.HI(tie_high_T28Y23), .LO(tie_low_T28Y23));
  sky130_fd_sc_hd__conb_1 conb_T28Y24 (.HI(tie_high_T28Y24), .LO(tie_low_T28Y24));
  sky130_fd_sc_hd__conb_1 conb_T28Y25 (.HI(tie_high_T28Y25), .LO(tie_low_T28Y25));
  sky130_fd_sc_hd__conb_1 conb_T28Y26 (.HI(tie_high_T28Y26), .LO(tie_low_T28Y26));
  sky130_fd_sc_hd__conb_1 conb_T28Y27 (.HI(tie_high_T28Y27), .LO(tie_low_T28Y27));
  sky130_fd_sc_hd__conb_1 conb_T28Y28 (.HI(tie_high_T28Y28), .LO(tie_low_T28Y28));
  sky130_fd_sc_hd__conb_1 conb_T28Y29 (.HI(tie_high_T28Y29), .LO(tie_low_T28Y29));
  sky130_fd_sc_hd__conb_1 conb_T28Y3 (.HI(tie_high_T28Y3), .LO(tie_low_T28Y3));
  sky130_fd_sc_hd__conb_1 conb_T28Y30 (.HI(tie_high_T28Y30), .LO(tie_low_T28Y30));
  sky130_fd_sc_hd__conb_1 conb_T28Y31 (.HI(tie_high_T28Y31), .LO(tie_low_T28Y31));
  sky130_fd_sc_hd__conb_1 conb_T28Y32 (.HI(tie_high_T28Y32), .LO(tie_low_T28Y32));
  sky130_fd_sc_hd__conb_1 conb_T28Y33 (.HI(tie_high_T28Y33), .LO(tie_low_T28Y33));
  sky130_fd_sc_hd__conb_1 conb_T28Y34 (.HI(tie_high_T28Y34), .LO(tie_low_T28Y34));
  sky130_fd_sc_hd__conb_1 conb_T28Y35 (.HI(tie_high_T28Y35), .LO(tie_low_T28Y35));
  sky130_fd_sc_hd__conb_1 conb_T28Y36 (.HI(tie_high_T28Y36), .LO(tie_low_T28Y36));
  sky130_fd_sc_hd__conb_1 conb_T28Y37 (.HI(tie_high_T28Y37), .LO(tie_low_T28Y37));
  sky130_fd_sc_hd__conb_1 conb_T28Y38 (.HI(tie_high_T28Y38), .LO(tie_low_T28Y38));
  sky130_fd_sc_hd__conb_1 conb_T28Y39 (.HI(tie_high_T28Y39), .LO(tie_low_T28Y39));
  sky130_fd_sc_hd__conb_1 conb_T28Y4 (.HI(tie_high_T28Y4), .LO(tie_low_T28Y4));
  sky130_fd_sc_hd__conb_1 conb_T28Y40 (.HI(tie_high_T28Y40), .LO(tie_low_T28Y40));
  sky130_fd_sc_hd__conb_1 conb_T28Y41 (.HI(tie_high_T28Y41), .LO(tie_low_T28Y41));
  sky130_fd_sc_hd__conb_1 conb_T28Y42 (.HI(tie_high_T28Y42), .LO(tie_low_T28Y42));
  sky130_fd_sc_hd__conb_1 conb_T28Y43 (.HI(tie_high_T28Y43), .LO(tie_low_T28Y43));
  sky130_fd_sc_hd__conb_1 conb_T28Y44 (.HI(tie_high_T28Y44), .LO(tie_low_T28Y44));
  sky130_fd_sc_hd__conb_1 conb_T28Y45 (.HI(tie_high_T28Y45), .LO(tie_low_T28Y45));
  sky130_fd_sc_hd__conb_1 conb_T28Y46 (.HI(tie_high_T28Y46), .LO(tie_low_T28Y46));
  sky130_fd_sc_hd__conb_1 conb_T28Y47 (.HI(tie_high_T28Y47), .LO(tie_low_T28Y47));
  sky130_fd_sc_hd__conb_1 conb_T28Y48 (.HI(tie_high_T28Y48), .LO(tie_low_T28Y48));
  sky130_fd_sc_hd__conb_1 conb_T28Y49 (.HI(tie_high_T28Y49), .LO(tie_low_T28Y49));
  sky130_fd_sc_hd__conb_1 conb_T28Y5 (.HI(tie_high_T28Y5), .LO(tie_low_T28Y5));
  sky130_fd_sc_hd__conb_1 conb_T28Y50 (.HI(tie_high_T28Y50), .LO(tie_low_T28Y50));
  sky130_fd_sc_hd__conb_1 conb_T28Y51 (.HI(tie_high_T28Y51), .LO(tie_low_T28Y51));
  sky130_fd_sc_hd__conb_1 conb_T28Y52 (.HI(tie_high_T28Y52), .LO(tie_low_T28Y52));
  sky130_fd_sc_hd__conb_1 conb_T28Y53 (.HI(tie_high_T28Y53), .LO(tie_low_T28Y53));
  sky130_fd_sc_hd__conb_1 conb_T28Y54 (.HI(tie_high_T28Y54), .LO(tie_low_T28Y54));
  sky130_fd_sc_hd__conb_1 conb_T28Y55 (.HI(tie_high_T28Y55), .LO(tie_low_T28Y55));
  sky130_fd_sc_hd__conb_1 conb_T28Y56 (.HI(tie_high_T28Y56), .LO(tie_low_T28Y56));
  sky130_fd_sc_hd__conb_1 conb_T28Y57 (.HI(tie_high_T28Y57), .LO(tie_low_T28Y57));
  sky130_fd_sc_hd__conb_1 conb_T28Y58 (.HI(tie_high_T28Y58), .LO(tie_low_T28Y58));
  sky130_fd_sc_hd__conb_1 conb_T28Y59 (.HI(tie_high_T28Y59), .LO(tie_low_T28Y59));
  sky130_fd_sc_hd__conb_1 conb_T28Y6 (.HI(tie_high_T28Y6), .LO(tie_low_T28Y6));
  sky130_fd_sc_hd__conb_1 conb_T28Y60 (.HI(tie_high_T28Y60), .LO(tie_low_T28Y60));
  sky130_fd_sc_hd__conb_1 conb_T28Y61 (.HI(tie_high_T28Y61), .LO(tie_low_T28Y61));
  sky130_fd_sc_hd__conb_1 conb_T28Y62 (.HI(tie_high_T28Y62), .LO(tie_low_T28Y62));
  sky130_fd_sc_hd__conb_1 conb_T28Y63 (.HI(tie_high_T28Y63), .LO(tie_low_T28Y63));
  sky130_fd_sc_hd__conb_1 conb_T28Y64 (.HI(tie_high_T28Y64), .LO(tie_low_T28Y64));
  sky130_fd_sc_hd__conb_1 conb_T28Y65 (.HI(tie_high_T28Y65), .LO(tie_low_T28Y65));
  sky130_fd_sc_hd__conb_1 conb_T28Y66 (.HI(tie_high_T28Y66), .LO(tie_low_T28Y66));
  sky130_fd_sc_hd__conb_1 conb_T28Y67 (.HI(tie_high_T28Y67), .LO(tie_low_T28Y67));
  sky130_fd_sc_hd__conb_1 conb_T28Y68 (.HI(tie_high_T28Y68), .LO(tie_low_T28Y68));
  sky130_fd_sc_hd__conb_1 conb_T28Y69 (.HI(tie_high_T28Y69), .LO(tie_low_T28Y69));
  sky130_fd_sc_hd__conb_1 conb_T28Y7 (.HI(tie_high_T28Y7), .LO(tie_low_T28Y7));
  sky130_fd_sc_hd__conb_1 conb_T28Y70 (.HI(tie_high_T28Y70), .LO(tie_low_T28Y70));
  sky130_fd_sc_hd__conb_1 conb_T28Y71 (.HI(tie_high_T28Y71), .LO(tie_low_T28Y71));
  sky130_fd_sc_hd__conb_1 conb_T28Y72 (.HI(tie_high_T28Y72), .LO(tie_low_T28Y72));
  sky130_fd_sc_hd__conb_1 conb_T28Y73 (.HI(tie_high_T28Y73), .LO(tie_low_T28Y73));
  sky130_fd_sc_hd__conb_1 conb_T28Y74 (.HI(tie_high_T28Y74), .LO(tie_low_T28Y74));
  sky130_fd_sc_hd__conb_1 conb_T28Y75 (.HI(tie_high_T28Y75), .LO(tie_low_T28Y75));
  sky130_fd_sc_hd__conb_1 conb_T28Y76 (.HI(tie_high_T28Y76), .LO(tie_low_T28Y76));
  sky130_fd_sc_hd__conb_1 conb_T28Y77 (.HI(tie_high_T28Y77), .LO(tie_low_T28Y77));
  sky130_fd_sc_hd__conb_1 conb_T28Y78 (.HI(tie_high_T28Y78), .LO(tie_low_T28Y78));
  sky130_fd_sc_hd__conb_1 conb_T28Y79 (.HI(tie_high_T28Y79), .LO(tie_low_T28Y79));
  sky130_fd_sc_hd__conb_1 conb_T28Y8 (.HI(tie_high_T28Y8), .LO(tie_low_T28Y8));
  sky130_fd_sc_hd__conb_1 conb_T28Y80 (.HI(tie_high_T28Y80), .LO(tie_low_T28Y80));
  sky130_fd_sc_hd__conb_1 conb_T28Y81 (.HI(tie_high_T28Y81), .LO(tie_low_T28Y81));
  sky130_fd_sc_hd__conb_1 conb_T28Y82 (.HI(tie_high_T28Y82), .LO(tie_low_T28Y82));
  sky130_fd_sc_hd__conb_1 conb_T28Y83 (.HI(tie_high_T28Y83), .LO(tie_low_T28Y83));
  sky130_fd_sc_hd__conb_1 conb_T28Y84 (.HI(tie_high_T28Y84), .LO(tie_low_T28Y84));
  sky130_fd_sc_hd__conb_1 conb_T28Y85 (.HI(tie_high_T28Y85), .LO(tie_low_T28Y85));
  sky130_fd_sc_hd__conb_1 conb_T28Y86 (.HI(tie_high_T28Y86), .LO(tie_low_T28Y86));
  sky130_fd_sc_hd__conb_1 conb_T28Y87 (.HI(tie_high_T28Y87), .LO(tie_low_T28Y87));
  sky130_fd_sc_hd__conb_1 conb_T28Y88 (.HI(tie_high_T28Y88), .LO(tie_low_T28Y88));
  sky130_fd_sc_hd__conb_1 conb_T28Y89 (.HI(tie_high_T28Y89), .LO(tie_low_T28Y89));
  sky130_fd_sc_hd__conb_1 conb_T28Y9 (.HI(tie_high_T28Y9), .LO(tie_low_T28Y9));
  sky130_fd_sc_hd__conb_1 conb_T29Y0 (.HI(tie_high_T29Y0), .LO(tie_low_T29Y0));
  sky130_fd_sc_hd__conb_1 conb_T29Y1 (.HI(tie_high_T29Y1), .LO(tie_low_T29Y1));
  sky130_fd_sc_hd__conb_1 conb_T29Y10 (.HI(tie_high_T29Y10), .LO(tie_low_T29Y10));
  sky130_fd_sc_hd__conb_1 conb_T29Y11 (.HI(tie_high_T29Y11), .LO(tie_low_T29Y11));
  sky130_fd_sc_hd__conb_1 conb_T29Y12 (.HI(tie_high_T29Y12), .LO(tie_low_T29Y12));
  sky130_fd_sc_hd__conb_1 conb_T29Y13 (.HI(tie_high_T29Y13), .LO(tie_low_T29Y13));
  sky130_fd_sc_hd__conb_1 conb_T29Y14 (.HI(tie_high_T29Y14), .LO(tie_low_T29Y14));
  sky130_fd_sc_hd__conb_1 conb_T29Y15 (.HI(tie_high_T29Y15), .LO(tie_low_T29Y15));
  sky130_fd_sc_hd__conb_1 conb_T29Y16 (.HI(tie_high_T29Y16), .LO(tie_low_T29Y16));
  sky130_fd_sc_hd__conb_1 conb_T29Y17 (.HI(tie_high_T29Y17), .LO(tie_low_T29Y17));
  sky130_fd_sc_hd__conb_1 conb_T29Y18 (.HI(tie_high_T29Y18), .LO(tie_low_T29Y18));
  sky130_fd_sc_hd__conb_1 conb_T29Y19 (.HI(tie_high_T29Y19), .LO(tie_low_T29Y19));
  sky130_fd_sc_hd__conb_1 conb_T29Y2 (.HI(tie_high_T29Y2), .LO(tie_low_T29Y2));
  sky130_fd_sc_hd__conb_1 conb_T29Y20 (.HI(tie_high_T29Y20), .LO(tie_low_T29Y20));
  sky130_fd_sc_hd__conb_1 conb_T29Y21 (.HI(tie_high_T29Y21), .LO(tie_low_T29Y21));
  sky130_fd_sc_hd__conb_1 conb_T29Y22 (.HI(tie_high_T29Y22), .LO(tie_low_T29Y22));
  sky130_fd_sc_hd__conb_1 conb_T29Y23 (.HI(tie_high_T29Y23), .LO(tie_low_T29Y23));
  sky130_fd_sc_hd__conb_1 conb_T29Y24 (.HI(tie_high_T29Y24), .LO(tie_low_T29Y24));
  sky130_fd_sc_hd__conb_1 conb_T29Y25 (.HI(tie_high_T29Y25), .LO(tie_low_T29Y25));
  sky130_fd_sc_hd__conb_1 conb_T29Y26 (.HI(tie_high_T29Y26), .LO(tie_low_T29Y26));
  sky130_fd_sc_hd__conb_1 conb_T29Y27 (.HI(tie_high_T29Y27), .LO(tie_low_T29Y27));
  sky130_fd_sc_hd__conb_1 conb_T29Y28 (.HI(tie_high_T29Y28), .LO(tie_low_T29Y28));
  sky130_fd_sc_hd__conb_1 conb_T29Y29 (.HI(tie_high_T29Y29), .LO(tie_low_T29Y29));
  sky130_fd_sc_hd__conb_1 conb_T29Y3 (.HI(tie_high_T29Y3), .LO(tie_low_T29Y3));
  sky130_fd_sc_hd__conb_1 conb_T29Y30 (.HI(tie_high_T29Y30), .LO(tie_low_T29Y30));
  sky130_fd_sc_hd__conb_1 conb_T29Y31 (.HI(tie_high_T29Y31), .LO(tie_low_T29Y31));
  sky130_fd_sc_hd__conb_1 conb_T29Y32 (.HI(tie_high_T29Y32), .LO(tie_low_T29Y32));
  sky130_fd_sc_hd__conb_1 conb_T29Y33 (.HI(tie_high_T29Y33), .LO(tie_low_T29Y33));
  sky130_fd_sc_hd__conb_1 conb_T29Y34 (.HI(tie_high_T29Y34), .LO(tie_low_T29Y34));
  sky130_fd_sc_hd__conb_1 conb_T29Y35 (.HI(tie_high_T29Y35), .LO(tie_low_T29Y35));
  sky130_fd_sc_hd__conb_1 conb_T29Y36 (.HI(tie_high_T29Y36), .LO(tie_low_T29Y36));
  sky130_fd_sc_hd__conb_1 conb_T29Y37 (.HI(tie_high_T29Y37), .LO(tie_low_T29Y37));
  sky130_fd_sc_hd__conb_1 conb_T29Y38 (.HI(tie_high_T29Y38), .LO(tie_low_T29Y38));
  sky130_fd_sc_hd__conb_1 conb_T29Y39 (.HI(tie_high_T29Y39), .LO(tie_low_T29Y39));
  sky130_fd_sc_hd__conb_1 conb_T29Y4 (.HI(tie_high_T29Y4), .LO(tie_low_T29Y4));
  sky130_fd_sc_hd__conb_1 conb_T29Y40 (.HI(tie_high_T29Y40), .LO(tie_low_T29Y40));
  sky130_fd_sc_hd__conb_1 conb_T29Y41 (.HI(tie_high_T29Y41), .LO(tie_low_T29Y41));
  sky130_fd_sc_hd__conb_1 conb_T29Y42 (.HI(tie_high_T29Y42), .LO(tie_low_T29Y42));
  sky130_fd_sc_hd__conb_1 conb_T29Y43 (.HI(tie_high_T29Y43), .LO(tie_low_T29Y43));
  sky130_fd_sc_hd__conb_1 conb_T29Y44 (.HI(tie_high_T29Y44), .LO(tie_low_T29Y44));
  sky130_fd_sc_hd__conb_1 conb_T29Y45 (.HI(tie_high_T29Y45), .LO(tie_low_T29Y45));
  sky130_fd_sc_hd__conb_1 conb_T29Y46 (.HI(tie_high_T29Y46), .LO(tie_low_T29Y46));
  sky130_fd_sc_hd__conb_1 conb_T29Y47 (.HI(tie_high_T29Y47), .LO(tie_low_T29Y47));
  sky130_fd_sc_hd__conb_1 conb_T29Y48 (.HI(tie_high_T29Y48), .LO(tie_low_T29Y48));
  sky130_fd_sc_hd__conb_1 conb_T29Y49 (.HI(tie_high_T29Y49), .LO(tie_low_T29Y49));
  sky130_fd_sc_hd__conb_1 conb_T29Y5 (.HI(tie_high_T29Y5), .LO(tie_low_T29Y5));
  sky130_fd_sc_hd__conb_1 conb_T29Y50 (.HI(tie_high_T29Y50), .LO(tie_low_T29Y50));
  sky130_fd_sc_hd__conb_1 conb_T29Y51 (.HI(tie_high_T29Y51), .LO(tie_low_T29Y51));
  sky130_fd_sc_hd__conb_1 conb_T29Y52 (.HI(tie_high_T29Y52), .LO(tie_low_T29Y52));
  sky130_fd_sc_hd__conb_1 conb_T29Y53 (.HI(tie_high_T29Y53), .LO(tie_low_T29Y53));
  sky130_fd_sc_hd__conb_1 conb_T29Y54 (.HI(tie_high_T29Y54), .LO(tie_low_T29Y54));
  sky130_fd_sc_hd__conb_1 conb_T29Y55 (.HI(tie_high_T29Y55), .LO(tie_low_T29Y55));
  sky130_fd_sc_hd__conb_1 conb_T29Y56 (.HI(tie_high_T29Y56), .LO(tie_low_T29Y56));
  sky130_fd_sc_hd__conb_1 conb_T29Y57 (.HI(tie_high_T29Y57), .LO(tie_low_T29Y57));
  sky130_fd_sc_hd__conb_1 conb_T29Y58 (.HI(tie_high_T29Y58), .LO(tie_low_T29Y58));
  sky130_fd_sc_hd__conb_1 conb_T29Y59 (.HI(tie_high_T29Y59), .LO(tie_low_T29Y59));
  sky130_fd_sc_hd__conb_1 conb_T29Y6 (.HI(tie_high_T29Y6), .LO(tie_low_T29Y6));
  sky130_fd_sc_hd__conb_1 conb_T29Y60 (.HI(tie_high_T29Y60), .LO(tie_low_T29Y60));
  sky130_fd_sc_hd__conb_1 conb_T29Y61 (.HI(tie_high_T29Y61), .LO(tie_low_T29Y61));
  sky130_fd_sc_hd__conb_1 conb_T29Y62 (.HI(tie_high_T29Y62), .LO(tie_low_T29Y62));
  sky130_fd_sc_hd__conb_1 conb_T29Y63 (.HI(tie_high_T29Y63), .LO(tie_low_T29Y63));
  sky130_fd_sc_hd__conb_1 conb_T29Y64 (.HI(tie_high_T29Y64), .LO(tie_low_T29Y64));
  sky130_fd_sc_hd__conb_1 conb_T29Y65 (.HI(tie_high_T29Y65), .LO(tie_low_T29Y65));
  sky130_fd_sc_hd__conb_1 conb_T29Y66 (.HI(tie_high_T29Y66), .LO(tie_low_T29Y66));
  sky130_fd_sc_hd__conb_1 conb_T29Y67 (.HI(tie_high_T29Y67), .LO(tie_low_T29Y67));
  sky130_fd_sc_hd__conb_1 conb_T29Y68 (.HI(tie_high_T29Y68), .LO(tie_low_T29Y68));
  sky130_fd_sc_hd__conb_1 conb_T29Y69 (.HI(tie_high_T29Y69), .LO(tie_low_T29Y69));
  sky130_fd_sc_hd__conb_1 conb_T29Y7 (.HI(tie_high_T29Y7), .LO(tie_low_T29Y7));
  sky130_fd_sc_hd__conb_1 conb_T29Y70 (.HI(tie_high_T29Y70), .LO(tie_low_T29Y70));
  sky130_fd_sc_hd__conb_1 conb_T29Y71 (.HI(tie_high_T29Y71), .LO(tie_low_T29Y71));
  sky130_fd_sc_hd__conb_1 conb_T29Y72 (.HI(tie_high_T29Y72), .LO(tie_low_T29Y72));
  sky130_fd_sc_hd__conb_1 conb_T29Y73 (.HI(tie_high_T29Y73), .LO(tie_low_T29Y73));
  sky130_fd_sc_hd__conb_1 conb_T29Y74 (.HI(tie_high_T29Y74), .LO(tie_low_T29Y74));
  sky130_fd_sc_hd__conb_1 conb_T29Y75 (.HI(tie_high_T29Y75), .LO(tie_low_T29Y75));
  sky130_fd_sc_hd__conb_1 conb_T29Y76 (.HI(tie_high_T29Y76), .LO(tie_low_T29Y76));
  sky130_fd_sc_hd__conb_1 conb_T29Y77 (.HI(tie_high_T29Y77), .LO(tie_low_T29Y77));
  sky130_fd_sc_hd__conb_1 conb_T29Y78 (.HI(tie_high_T29Y78), .LO(tie_low_T29Y78));
  sky130_fd_sc_hd__conb_1 conb_T29Y79 (.HI(tie_high_T29Y79), .LO(tie_low_T29Y79));
  sky130_fd_sc_hd__conb_1 conb_T29Y8 (.HI(tie_high_T29Y8), .LO(tie_low_T29Y8));
  sky130_fd_sc_hd__conb_1 conb_T29Y80 (.HI(tie_high_T29Y80), .LO(tie_low_T29Y80));
  sky130_fd_sc_hd__conb_1 conb_T29Y81 (.HI(tie_high_T29Y81), .LO(tie_low_T29Y81));
  sky130_fd_sc_hd__conb_1 conb_T29Y82 (.HI(tie_high_T29Y82), .LO(tie_low_T29Y82));
  sky130_fd_sc_hd__conb_1 conb_T29Y83 (.HI(tie_high_T29Y83), .LO(tie_low_T29Y83));
  sky130_fd_sc_hd__conb_1 conb_T29Y84 (.HI(tie_high_T29Y84), .LO(tie_low_T29Y84));
  sky130_fd_sc_hd__conb_1 conb_T29Y85 (.HI(tie_high_T29Y85), .LO(tie_low_T29Y85));
  sky130_fd_sc_hd__conb_1 conb_T29Y86 (.HI(tie_high_T29Y86), .LO(tie_low_T29Y86));
  sky130_fd_sc_hd__conb_1 conb_T29Y87 (.HI(tie_high_T29Y87), .LO(tie_low_T29Y87));
  sky130_fd_sc_hd__conb_1 conb_T29Y88 (.HI(tie_high_T29Y88), .LO(tie_low_T29Y88));
  sky130_fd_sc_hd__conb_1 conb_T29Y89 (.HI(tie_high_T29Y89), .LO(tie_low_T29Y89));
  sky130_fd_sc_hd__conb_1 conb_T29Y9 (.HI(tie_high_T29Y9), .LO(tie_low_T29Y9));
  sky130_fd_sc_hd__conb_1 conb_T2Y0 (.HI(tie_high_T2Y0), .LO(tie_low_T2Y0));
  sky130_fd_sc_hd__conb_1 conb_T2Y1 (.HI(tie_high_T2Y1), .LO(tie_low_T2Y1));
  sky130_fd_sc_hd__conb_1 conb_T2Y10 (.HI(tie_high_T2Y10), .LO(tie_low_T2Y10));
  sky130_fd_sc_hd__conb_1 conb_T2Y11 (.HI(tie_high_T2Y11), .LO(tie_low_T2Y11));
  sky130_fd_sc_hd__conb_1 conb_T2Y12 (.HI(tie_high_T2Y12), .LO(tie_low_T2Y12));
  sky130_fd_sc_hd__conb_1 conb_T2Y13 (.HI(tie_high_T2Y13), .LO(tie_low_T2Y13));
  sky130_fd_sc_hd__conb_1 conb_T2Y14 (.HI(tie_high_T2Y14), .LO(tie_low_T2Y14));
  sky130_fd_sc_hd__conb_1 conb_T2Y15 (.HI(tie_high_T2Y15), .LO(tie_low_T2Y15));
  sky130_fd_sc_hd__conb_1 conb_T2Y16 (.HI(tie_high_T2Y16), .LO(tie_low_T2Y16));
  sky130_fd_sc_hd__conb_1 conb_T2Y17 (.HI(tie_high_T2Y17), .LO(tie_low_T2Y17));
  sky130_fd_sc_hd__conb_1 conb_T2Y18 (.HI(tie_high_T2Y18), .LO(tie_low_T2Y18));
  sky130_fd_sc_hd__conb_1 conb_T2Y19 (.HI(tie_high_T2Y19), .LO(tie_low_T2Y19));
  sky130_fd_sc_hd__conb_1 conb_T2Y2 (.HI(tie_high_T2Y2), .LO(tie_low_T2Y2));
  sky130_fd_sc_hd__conb_1 conb_T2Y20 (.HI(tie_high_T2Y20), .LO(tie_low_T2Y20));
  sky130_fd_sc_hd__conb_1 conb_T2Y21 (.HI(tie_high_T2Y21), .LO(tie_low_T2Y21));
  sky130_fd_sc_hd__conb_1 conb_T2Y22 (.HI(tie_high_T2Y22), .LO(tie_low_T2Y22));
  sky130_fd_sc_hd__conb_1 conb_T2Y23 (.HI(tie_high_T2Y23), .LO(tie_low_T2Y23));
  sky130_fd_sc_hd__conb_1 conb_T2Y24 (.HI(tie_high_T2Y24), .LO(tie_low_T2Y24));
  sky130_fd_sc_hd__conb_1 conb_T2Y25 (.HI(tie_high_T2Y25), .LO(tie_low_T2Y25));
  sky130_fd_sc_hd__conb_1 conb_T2Y26 (.HI(tie_high_T2Y26), .LO(tie_low_T2Y26));
  sky130_fd_sc_hd__conb_1 conb_T2Y27 (.HI(tie_high_T2Y27), .LO(tie_low_T2Y27));
  sky130_fd_sc_hd__conb_1 conb_T2Y28 (.HI(tie_high_T2Y28), .LO(tie_low_T2Y28));
  sky130_fd_sc_hd__conb_1 conb_T2Y29 (.HI(tie_high_T2Y29), .LO(tie_low_T2Y29));
  sky130_fd_sc_hd__conb_1 conb_T2Y3 (.HI(tie_high_T2Y3), .LO(tie_low_T2Y3));
  sky130_fd_sc_hd__conb_1 conb_T2Y30 (.HI(tie_high_T2Y30), .LO(tie_low_T2Y30));
  sky130_fd_sc_hd__conb_1 conb_T2Y31 (.HI(tie_high_T2Y31), .LO(tie_low_T2Y31));
  sky130_fd_sc_hd__conb_1 conb_T2Y32 (.HI(tie_high_T2Y32), .LO(tie_low_T2Y32));
  sky130_fd_sc_hd__conb_1 conb_T2Y33 (.HI(tie_high_T2Y33), .LO(tie_low_T2Y33));
  sky130_fd_sc_hd__conb_1 conb_T2Y34 (.HI(tie_high_T2Y34), .LO(tie_low_T2Y34));
  sky130_fd_sc_hd__conb_1 conb_T2Y35 (.HI(tie_high_T2Y35), .LO(tie_low_T2Y35));
  sky130_fd_sc_hd__conb_1 conb_T2Y36 (.HI(tie_high_T2Y36), .LO(tie_low_T2Y36));
  sky130_fd_sc_hd__conb_1 conb_T2Y37 (.HI(tie_high_T2Y37), .LO(tie_low_T2Y37));
  sky130_fd_sc_hd__conb_1 conb_T2Y38 (.HI(tie_high_T2Y38), .LO(tie_low_T2Y38));
  sky130_fd_sc_hd__conb_1 conb_T2Y39 (.HI(tie_high_T2Y39), .LO(tie_low_T2Y39));
  sky130_fd_sc_hd__conb_1 conb_T2Y4 (.HI(tie_high_T2Y4), .LO(tie_low_T2Y4));
  sky130_fd_sc_hd__conb_1 conb_T2Y40 (.HI(tie_high_T2Y40), .LO(tie_low_T2Y40));
  sky130_fd_sc_hd__conb_1 conb_T2Y41 (.HI(tie_high_T2Y41), .LO(tie_low_T2Y41));
  sky130_fd_sc_hd__conb_1 conb_T2Y42 (.HI(tie_high_T2Y42), .LO(tie_low_T2Y42));
  sky130_fd_sc_hd__conb_1 conb_T2Y43 (.HI(tie_high_T2Y43), .LO(tie_low_T2Y43));
  sky130_fd_sc_hd__conb_1 conb_T2Y44 (.HI(tie_high_T2Y44), .LO(tie_low_T2Y44));
  sky130_fd_sc_hd__conb_1 conb_T2Y45 (.HI(tie_high_T2Y45), .LO(tie_low_T2Y45));
  sky130_fd_sc_hd__conb_1 conb_T2Y46 (.HI(tie_high_T2Y46), .LO(tie_low_T2Y46));
  sky130_fd_sc_hd__conb_1 conb_T2Y47 (.HI(tie_high_T2Y47), .LO(tie_low_T2Y47));
  sky130_fd_sc_hd__conb_1 conb_T2Y48 (.HI(tie_high_T2Y48), .LO(tie_low_T2Y48));
  sky130_fd_sc_hd__conb_1 conb_T2Y49 (.HI(tie_high_T2Y49), .LO(tie_low_T2Y49));
  sky130_fd_sc_hd__conb_1 conb_T2Y5 (.HI(tie_high_T2Y5), .LO(tie_low_T2Y5));
  sky130_fd_sc_hd__conb_1 conb_T2Y50 (.HI(tie_high_T2Y50), .LO(tie_low_T2Y50));
  sky130_fd_sc_hd__conb_1 conb_T2Y51 (.HI(tie_high_T2Y51), .LO(tie_low_T2Y51));
  sky130_fd_sc_hd__conb_1 conb_T2Y52 (.HI(tie_high_T2Y52), .LO(tie_low_T2Y52));
  sky130_fd_sc_hd__conb_1 conb_T2Y53 (.HI(tie_high_T2Y53), .LO(tie_low_T2Y53));
  sky130_fd_sc_hd__conb_1 conb_T2Y54 (.HI(tie_high_T2Y54), .LO(tie_low_T2Y54));
  sky130_fd_sc_hd__conb_1 conb_T2Y55 (.HI(tie_high_T2Y55), .LO(tie_low_T2Y55));
  sky130_fd_sc_hd__conb_1 conb_T2Y56 (.HI(tie_high_T2Y56), .LO(tie_low_T2Y56));
  sky130_fd_sc_hd__conb_1 conb_T2Y57 (.HI(tie_high_T2Y57), .LO(tie_low_T2Y57));
  sky130_fd_sc_hd__conb_1 conb_T2Y58 (.HI(tie_high_T2Y58), .LO(tie_low_T2Y58));
  sky130_fd_sc_hd__conb_1 conb_T2Y59 (.HI(tie_high_T2Y59), .LO(tie_low_T2Y59));
  sky130_fd_sc_hd__conb_1 conb_T2Y6 (.HI(tie_high_T2Y6), .LO(tie_low_T2Y6));
  sky130_fd_sc_hd__conb_1 conb_T2Y60 (.HI(tie_high_T2Y60), .LO(tie_low_T2Y60));
  sky130_fd_sc_hd__conb_1 conb_T2Y61 (.HI(tie_high_T2Y61), .LO(tie_low_T2Y61));
  sky130_fd_sc_hd__conb_1 conb_T2Y62 (.HI(tie_high_T2Y62), .LO(tie_low_T2Y62));
  sky130_fd_sc_hd__conb_1 conb_T2Y63 (.HI(tie_high_T2Y63), .LO(tie_low_T2Y63));
  sky130_fd_sc_hd__conb_1 conb_T2Y64 (.HI(tie_high_T2Y64), .LO(tie_low_T2Y64));
  sky130_fd_sc_hd__conb_1 conb_T2Y65 (.HI(tie_high_T2Y65), .LO(tie_low_T2Y65));
  sky130_fd_sc_hd__conb_1 conb_T2Y66 (.HI(tie_high_T2Y66), .LO(tie_low_T2Y66));
  sky130_fd_sc_hd__conb_1 conb_T2Y67 (.HI(tie_high_T2Y67), .LO(tie_low_T2Y67));
  sky130_fd_sc_hd__conb_1 conb_T2Y68 (.HI(tie_high_T2Y68), .LO(tie_low_T2Y68));
  sky130_fd_sc_hd__conb_1 conb_T2Y69 (.HI(tie_high_T2Y69), .LO(tie_low_T2Y69));
  sky130_fd_sc_hd__conb_1 conb_T2Y7 (.HI(tie_high_T2Y7), .LO(tie_low_T2Y7));
  sky130_fd_sc_hd__conb_1 conb_T2Y70 (.HI(tie_high_T2Y70), .LO(tie_low_T2Y70));
  sky130_fd_sc_hd__conb_1 conb_T2Y71 (.HI(tie_high_T2Y71), .LO(tie_low_T2Y71));
  sky130_fd_sc_hd__conb_1 conb_T2Y72 (.HI(tie_high_T2Y72), .LO(tie_low_T2Y72));
  sky130_fd_sc_hd__conb_1 conb_T2Y73 (.HI(tie_high_T2Y73), .LO(tie_low_T2Y73));
  sky130_fd_sc_hd__conb_1 conb_T2Y74 (.HI(tie_high_T2Y74), .LO(tie_low_T2Y74));
  sky130_fd_sc_hd__conb_1 conb_T2Y75 (.HI(tie_high_T2Y75), .LO(tie_low_T2Y75));
  sky130_fd_sc_hd__conb_1 conb_T2Y76 (.HI(tie_high_T2Y76), .LO(tie_low_T2Y76));
  sky130_fd_sc_hd__conb_1 conb_T2Y77 (.HI(tie_high_T2Y77), .LO(tie_low_T2Y77));
  sky130_fd_sc_hd__conb_1 conb_T2Y78 (.HI(tie_high_T2Y78), .LO(tie_low_T2Y78));
  sky130_fd_sc_hd__conb_1 conb_T2Y79 (.HI(tie_high_T2Y79), .LO(tie_low_T2Y79));
  sky130_fd_sc_hd__conb_1 conb_T2Y8 (.HI(tie_high_T2Y8), .LO(tie_low_T2Y8));
  sky130_fd_sc_hd__conb_1 conb_T2Y80 (.HI(tie_high_T2Y80), .LO(tie_low_T2Y80));
  sky130_fd_sc_hd__conb_1 conb_T2Y81 (.HI(tie_high_T2Y81), .LO(tie_low_T2Y81));
  sky130_fd_sc_hd__conb_1 conb_T2Y82 (.HI(tie_high_T2Y82), .LO(tie_low_T2Y82));
  sky130_fd_sc_hd__conb_1 conb_T2Y83 (.HI(tie_high_T2Y83), .LO(tie_low_T2Y83));
  sky130_fd_sc_hd__conb_1 conb_T2Y84 (.HI(tie_high_T2Y84), .LO(tie_low_T2Y84));
  sky130_fd_sc_hd__conb_1 conb_T2Y85 (.HI(tie_high_T2Y85), .LO(tie_low_T2Y85));
  sky130_fd_sc_hd__conb_1 conb_T2Y86 (.HI(tie_high_T2Y86), .LO(tie_low_T2Y86));
  sky130_fd_sc_hd__conb_1 conb_T2Y87 (.HI(tie_high_T2Y87), .LO(tie_low_T2Y87));
  sky130_fd_sc_hd__conb_1 conb_T2Y88 (.HI(tie_high_T2Y88), .LO(tie_low_T2Y88));
  sky130_fd_sc_hd__conb_1 conb_T2Y89 (.HI(tie_high_T2Y89), .LO(tie_low_T2Y89));
  sky130_fd_sc_hd__conb_1 conb_T2Y9 (.HI(tie_high_T2Y9), .LO(tie_low_T2Y9));
  sky130_fd_sc_hd__conb_1 conb_T30Y0 (.HI(tie_high_T30Y0), .LO(tie_low_T30Y0));
  sky130_fd_sc_hd__conb_1 conb_T30Y1 (.HI(tie_high_T30Y1), .LO(tie_low_T30Y1));
  sky130_fd_sc_hd__conb_1 conb_T30Y10 (.HI(tie_high_T30Y10), .LO(tie_low_T30Y10));
  sky130_fd_sc_hd__conb_1 conb_T30Y11 (.HI(tie_high_T30Y11), .LO(tie_low_T30Y11));
  sky130_fd_sc_hd__conb_1 conb_T30Y12 (.HI(tie_high_T30Y12), .LO(tie_low_T30Y12));
  sky130_fd_sc_hd__conb_1 conb_T30Y13 (.HI(tie_high_T30Y13), .LO(tie_low_T30Y13));
  sky130_fd_sc_hd__conb_1 conb_T30Y14 (.HI(tie_high_T30Y14), .LO(tie_low_T30Y14));
  sky130_fd_sc_hd__conb_1 conb_T30Y15 (.HI(tie_high_T30Y15), .LO(tie_low_T30Y15));
  sky130_fd_sc_hd__conb_1 conb_T30Y16 (.HI(tie_high_T30Y16), .LO(tie_low_T30Y16));
  sky130_fd_sc_hd__conb_1 conb_T30Y17 (.HI(tie_high_T30Y17), .LO(tie_low_T30Y17));
  sky130_fd_sc_hd__conb_1 conb_T30Y18 (.HI(tie_high_T30Y18), .LO(tie_low_T30Y18));
  sky130_fd_sc_hd__conb_1 conb_T30Y19 (.HI(tie_high_T30Y19), .LO(tie_low_T30Y19));
  sky130_fd_sc_hd__conb_1 conb_T30Y2 (.HI(tie_high_T30Y2), .LO(tie_low_T30Y2));
  sky130_fd_sc_hd__conb_1 conb_T30Y20 (.HI(tie_high_T30Y20), .LO(tie_low_T30Y20));
  sky130_fd_sc_hd__conb_1 conb_T30Y21 (.HI(tie_high_T30Y21), .LO(tie_low_T30Y21));
  sky130_fd_sc_hd__conb_1 conb_T30Y22 (.HI(tie_high_T30Y22), .LO(tie_low_T30Y22));
  sky130_fd_sc_hd__conb_1 conb_T30Y23 (.HI(tie_high_T30Y23), .LO(tie_low_T30Y23));
  sky130_fd_sc_hd__conb_1 conb_T30Y24 (.HI(tie_high_T30Y24), .LO(tie_low_T30Y24));
  sky130_fd_sc_hd__conb_1 conb_T30Y25 (.HI(tie_high_T30Y25), .LO(tie_low_T30Y25));
  sky130_fd_sc_hd__conb_1 conb_T30Y26 (.HI(tie_high_T30Y26), .LO(tie_low_T30Y26));
  sky130_fd_sc_hd__conb_1 conb_T30Y27 (.HI(tie_high_T30Y27), .LO(tie_low_T30Y27));
  sky130_fd_sc_hd__conb_1 conb_T30Y28 (.HI(tie_high_T30Y28), .LO(tie_low_T30Y28));
  sky130_fd_sc_hd__conb_1 conb_T30Y29 (.HI(tie_high_T30Y29), .LO(tie_low_T30Y29));
  sky130_fd_sc_hd__conb_1 conb_T30Y3 (.HI(tie_high_T30Y3), .LO(tie_low_T30Y3));
  sky130_fd_sc_hd__conb_1 conb_T30Y30 (.HI(tie_high_T30Y30), .LO(tie_low_T30Y30));
  sky130_fd_sc_hd__conb_1 conb_T30Y31 (.HI(tie_high_T30Y31), .LO(tie_low_T30Y31));
  sky130_fd_sc_hd__conb_1 conb_T30Y32 (.HI(tie_high_T30Y32), .LO(tie_low_T30Y32));
  sky130_fd_sc_hd__conb_1 conb_T30Y33 (.HI(tie_high_T30Y33), .LO(tie_low_T30Y33));
  sky130_fd_sc_hd__conb_1 conb_T30Y34 (.HI(tie_high_T30Y34), .LO(tie_low_T30Y34));
  sky130_fd_sc_hd__conb_1 conb_T30Y35 (.HI(tie_high_T30Y35), .LO(tie_low_T30Y35));
  sky130_fd_sc_hd__conb_1 conb_T30Y36 (.HI(tie_high_T30Y36), .LO(tie_low_T30Y36));
  sky130_fd_sc_hd__conb_1 conb_T30Y37 (.HI(tie_high_T30Y37), .LO(tie_low_T30Y37));
  sky130_fd_sc_hd__conb_1 conb_T30Y38 (.HI(tie_high_T30Y38), .LO(tie_low_T30Y38));
  sky130_fd_sc_hd__conb_1 conb_T30Y39 (.HI(tie_high_T30Y39), .LO(tie_low_T30Y39));
  sky130_fd_sc_hd__conb_1 conb_T30Y4 (.HI(tie_high_T30Y4), .LO(tie_low_T30Y4));
  sky130_fd_sc_hd__conb_1 conb_T30Y40 (.HI(tie_high_T30Y40), .LO(tie_low_T30Y40));
  sky130_fd_sc_hd__conb_1 conb_T30Y41 (.HI(tie_high_T30Y41), .LO(tie_low_T30Y41));
  sky130_fd_sc_hd__conb_1 conb_T30Y42 (.HI(tie_high_T30Y42), .LO(tie_low_T30Y42));
  sky130_fd_sc_hd__conb_1 conb_T30Y43 (.HI(tie_high_T30Y43), .LO(tie_low_T30Y43));
  sky130_fd_sc_hd__conb_1 conb_T30Y44 (.HI(tie_high_T30Y44), .LO(tie_low_T30Y44));
  sky130_fd_sc_hd__conb_1 conb_T30Y45 (.HI(tie_high_T30Y45), .LO(tie_low_T30Y45));
  sky130_fd_sc_hd__conb_1 conb_T30Y46 (.HI(tie_high_T30Y46), .LO(tie_low_T30Y46));
  sky130_fd_sc_hd__conb_1 conb_T30Y47 (.HI(tie_high_T30Y47), .LO(tie_low_T30Y47));
  sky130_fd_sc_hd__conb_1 conb_T30Y48 (.HI(tie_high_T30Y48), .LO(tie_low_T30Y48));
  sky130_fd_sc_hd__conb_1 conb_T30Y49 (.HI(tie_high_T30Y49), .LO(tie_low_T30Y49));
  sky130_fd_sc_hd__conb_1 conb_T30Y5 (.HI(tie_high_T30Y5), .LO(tie_low_T30Y5));
  sky130_fd_sc_hd__conb_1 conb_T30Y50 (.HI(tie_high_T30Y50), .LO(tie_low_T30Y50));
  sky130_fd_sc_hd__conb_1 conb_T30Y51 (.HI(tie_high_T30Y51), .LO(tie_low_T30Y51));
  sky130_fd_sc_hd__conb_1 conb_T30Y52 (.HI(tie_high_T30Y52), .LO(tie_low_T30Y52));
  sky130_fd_sc_hd__conb_1 conb_T30Y53 (.HI(tie_high_T30Y53), .LO(tie_low_T30Y53));
  sky130_fd_sc_hd__conb_1 conb_T30Y54 (.HI(tie_high_T30Y54), .LO(tie_low_T30Y54));
  sky130_fd_sc_hd__conb_1 conb_T30Y55 (.HI(tie_high_T30Y55), .LO(tie_low_T30Y55));
  sky130_fd_sc_hd__conb_1 conb_T30Y56 (.HI(tie_high_T30Y56), .LO(tie_low_T30Y56));
  sky130_fd_sc_hd__conb_1 conb_T30Y57 (.HI(tie_high_T30Y57), .LO(tie_low_T30Y57));
  sky130_fd_sc_hd__conb_1 conb_T30Y58 (.HI(tie_high_T30Y58), .LO(tie_low_T30Y58));
  sky130_fd_sc_hd__conb_1 conb_T30Y59 (.HI(tie_high_T30Y59), .LO(tie_low_T30Y59));
  sky130_fd_sc_hd__conb_1 conb_T30Y6 (.HI(tie_high_T30Y6), .LO(tie_low_T30Y6));
  sky130_fd_sc_hd__conb_1 conb_T30Y60 (.HI(tie_high_T30Y60), .LO(tie_low_T30Y60));
  sky130_fd_sc_hd__conb_1 conb_T30Y61 (.HI(tie_high_T30Y61), .LO(tie_low_T30Y61));
  sky130_fd_sc_hd__conb_1 conb_T30Y62 (.HI(tie_high_T30Y62), .LO(tie_low_T30Y62));
  sky130_fd_sc_hd__conb_1 conb_T30Y63 (.HI(tie_high_T30Y63), .LO(tie_low_T30Y63));
  sky130_fd_sc_hd__conb_1 conb_T30Y64 (.HI(tie_high_T30Y64), .LO(tie_low_T30Y64));
  sky130_fd_sc_hd__conb_1 conb_T30Y65 (.HI(tie_high_T30Y65), .LO(tie_low_T30Y65));
  sky130_fd_sc_hd__conb_1 conb_T30Y66 (.HI(tie_high_T30Y66), .LO(tie_low_T30Y66));
  sky130_fd_sc_hd__conb_1 conb_T30Y67 (.HI(tie_high_T30Y67), .LO(tie_low_T30Y67));
  sky130_fd_sc_hd__conb_1 conb_T30Y68 (.HI(tie_high_T30Y68), .LO(tie_low_T30Y68));
  sky130_fd_sc_hd__conb_1 conb_T30Y69 (.HI(tie_high_T30Y69), .LO(tie_low_T30Y69));
  sky130_fd_sc_hd__conb_1 conb_T30Y7 (.HI(tie_high_T30Y7), .LO(tie_low_T30Y7));
  sky130_fd_sc_hd__conb_1 conb_T30Y70 (.HI(tie_high_T30Y70), .LO(tie_low_T30Y70));
  sky130_fd_sc_hd__conb_1 conb_T30Y71 (.HI(tie_high_T30Y71), .LO(tie_low_T30Y71));
  sky130_fd_sc_hd__conb_1 conb_T30Y72 (.HI(tie_high_T30Y72), .LO(tie_low_T30Y72));
  sky130_fd_sc_hd__conb_1 conb_T30Y73 (.HI(tie_high_T30Y73), .LO(tie_low_T30Y73));
  sky130_fd_sc_hd__conb_1 conb_T30Y74 (.HI(tie_high_T30Y74), .LO(tie_low_T30Y74));
  sky130_fd_sc_hd__conb_1 conb_T30Y75 (.HI(tie_high_T30Y75), .LO(tie_low_T30Y75));
  sky130_fd_sc_hd__conb_1 conb_T30Y76 (.HI(tie_high_T30Y76), .LO(tie_low_T30Y76));
  sky130_fd_sc_hd__conb_1 conb_T30Y77 (.HI(tie_high_T30Y77), .LO(tie_low_T30Y77));
  sky130_fd_sc_hd__conb_1 conb_T30Y78 (.HI(tie_high_T30Y78), .LO(tie_low_T30Y78));
  sky130_fd_sc_hd__conb_1 conb_T30Y79 (.HI(tie_high_T30Y79), .LO(tie_low_T30Y79));
  sky130_fd_sc_hd__conb_1 conb_T30Y8 (.HI(tie_high_T30Y8), .LO(tie_low_T30Y8));
  sky130_fd_sc_hd__conb_1 conb_T30Y80 (.HI(tie_high_T30Y80), .LO(tie_low_T30Y80));
  sky130_fd_sc_hd__conb_1 conb_T30Y81 (.HI(tie_high_T30Y81), .LO(tie_low_T30Y81));
  sky130_fd_sc_hd__conb_1 conb_T30Y82 (.HI(tie_high_T30Y82), .LO(tie_low_T30Y82));
  sky130_fd_sc_hd__conb_1 conb_T30Y83 (.HI(tie_high_T30Y83), .LO(tie_low_T30Y83));
  sky130_fd_sc_hd__conb_1 conb_T30Y84 (.HI(tie_high_T30Y84), .LO(tie_low_T30Y84));
  sky130_fd_sc_hd__conb_1 conb_T30Y85 (.HI(tie_high_T30Y85), .LO(tie_low_T30Y85));
  sky130_fd_sc_hd__conb_1 conb_T30Y86 (.HI(tie_high_T30Y86), .LO(tie_low_T30Y86));
  sky130_fd_sc_hd__conb_1 conb_T30Y87 (.HI(tie_high_T30Y87), .LO(tie_low_T30Y87));
  sky130_fd_sc_hd__conb_1 conb_T30Y88 (.HI(tie_high_T30Y88), .LO(tie_low_T30Y88));
  sky130_fd_sc_hd__conb_1 conb_T30Y89 (.HI(tie_high_T30Y89), .LO(tie_low_T30Y89));
  sky130_fd_sc_hd__conb_1 conb_T30Y9 (.HI(tie_high_T30Y9), .LO(tie_low_T30Y9));
  sky130_fd_sc_hd__conb_1 conb_T31Y0 (.HI(tie_high_T31Y0), .LO(tie_low_T31Y0));
  sky130_fd_sc_hd__conb_1 conb_T31Y1 (.HI(tie_high_T31Y1), .LO(tie_low_T31Y1));
  sky130_fd_sc_hd__conb_1 conb_T31Y10 (.HI(tie_high_T31Y10), .LO(tie_low_T31Y10));
  sky130_fd_sc_hd__conb_1 conb_T31Y11 (.HI(tie_high_T31Y11), .LO(tie_low_T31Y11));
  sky130_fd_sc_hd__conb_1 conb_T31Y12 (.HI(tie_high_T31Y12), .LO(tie_low_T31Y12));
  sky130_fd_sc_hd__conb_1 conb_T31Y13 (.HI(tie_high_T31Y13), .LO(tie_low_T31Y13));
  sky130_fd_sc_hd__conb_1 conb_T31Y14 (.HI(tie_high_T31Y14), .LO(tie_low_T31Y14));
  sky130_fd_sc_hd__conb_1 conb_T31Y15 (.HI(tie_high_T31Y15), .LO(tie_low_T31Y15));
  sky130_fd_sc_hd__conb_1 conb_T31Y16 (.HI(tie_high_T31Y16), .LO(tie_low_T31Y16));
  sky130_fd_sc_hd__conb_1 conb_T31Y17 (.HI(tie_high_T31Y17), .LO(tie_low_T31Y17));
  sky130_fd_sc_hd__conb_1 conb_T31Y18 (.HI(tie_high_T31Y18), .LO(tie_low_T31Y18));
  sky130_fd_sc_hd__conb_1 conb_T31Y19 (.HI(tie_high_T31Y19), .LO(tie_low_T31Y19));
  sky130_fd_sc_hd__conb_1 conb_T31Y2 (.HI(tie_high_T31Y2), .LO(tie_low_T31Y2));
  sky130_fd_sc_hd__conb_1 conb_T31Y20 (.HI(tie_high_T31Y20), .LO(tie_low_T31Y20));
  sky130_fd_sc_hd__conb_1 conb_T31Y21 (.HI(tie_high_T31Y21), .LO(tie_low_T31Y21));
  sky130_fd_sc_hd__conb_1 conb_T31Y22 (.HI(tie_high_T31Y22), .LO(tie_low_T31Y22));
  sky130_fd_sc_hd__conb_1 conb_T31Y23 (.HI(tie_high_T31Y23), .LO(tie_low_T31Y23));
  sky130_fd_sc_hd__conb_1 conb_T31Y24 (.HI(tie_high_T31Y24), .LO(tie_low_T31Y24));
  sky130_fd_sc_hd__conb_1 conb_T31Y25 (.HI(tie_high_T31Y25), .LO(tie_low_T31Y25));
  sky130_fd_sc_hd__conb_1 conb_T31Y26 (.HI(tie_high_T31Y26), .LO(tie_low_T31Y26));
  sky130_fd_sc_hd__conb_1 conb_T31Y27 (.HI(tie_high_T31Y27), .LO(tie_low_T31Y27));
  sky130_fd_sc_hd__conb_1 conb_T31Y28 (.HI(tie_high_T31Y28), .LO(tie_low_T31Y28));
  sky130_fd_sc_hd__conb_1 conb_T31Y29 (.HI(tie_high_T31Y29), .LO(tie_low_T31Y29));
  sky130_fd_sc_hd__conb_1 conb_T31Y3 (.HI(tie_high_T31Y3), .LO(tie_low_T31Y3));
  sky130_fd_sc_hd__conb_1 conb_T31Y30 (.HI(tie_high_T31Y30), .LO(tie_low_T31Y30));
  sky130_fd_sc_hd__conb_1 conb_T31Y31 (.HI(tie_high_T31Y31), .LO(tie_low_T31Y31));
  sky130_fd_sc_hd__conb_1 conb_T31Y32 (.HI(tie_high_T31Y32), .LO(tie_low_T31Y32));
  sky130_fd_sc_hd__conb_1 conb_T31Y33 (.HI(tie_high_T31Y33), .LO(tie_low_T31Y33));
  sky130_fd_sc_hd__conb_1 conb_T31Y34 (.HI(tie_high_T31Y34), .LO(tie_low_T31Y34));
  sky130_fd_sc_hd__conb_1 conb_T31Y35 (.HI(tie_high_T31Y35), .LO(tie_low_T31Y35));
  sky130_fd_sc_hd__conb_1 conb_T31Y36 (.HI(tie_high_T31Y36), .LO(tie_low_T31Y36));
  sky130_fd_sc_hd__conb_1 conb_T31Y37 (.HI(tie_high_T31Y37), .LO(tie_low_T31Y37));
  sky130_fd_sc_hd__conb_1 conb_T31Y38 (.HI(tie_high_T31Y38), .LO(tie_low_T31Y38));
  sky130_fd_sc_hd__conb_1 conb_T31Y39 (.HI(tie_high_T31Y39), .LO(tie_low_T31Y39));
  sky130_fd_sc_hd__conb_1 conb_T31Y4 (.HI(tie_high_T31Y4), .LO(tie_low_T31Y4));
  sky130_fd_sc_hd__conb_1 conb_T31Y40 (.HI(tie_high_T31Y40), .LO(tie_low_T31Y40));
  sky130_fd_sc_hd__conb_1 conb_T31Y41 (.HI(tie_high_T31Y41), .LO(tie_low_T31Y41));
  sky130_fd_sc_hd__conb_1 conb_T31Y42 (.HI(tie_high_T31Y42), .LO(tie_low_T31Y42));
  sky130_fd_sc_hd__conb_1 conb_T31Y43 (.HI(tie_high_T31Y43), .LO(tie_low_T31Y43));
  sky130_fd_sc_hd__conb_1 conb_T31Y44 (.HI(tie_high_T31Y44), .LO(tie_low_T31Y44));
  sky130_fd_sc_hd__conb_1 conb_T31Y45 (.HI(tie_high_T31Y45), .LO(tie_low_T31Y45));
  sky130_fd_sc_hd__conb_1 conb_T31Y46 (.HI(tie_high_T31Y46), .LO(tie_low_T31Y46));
  sky130_fd_sc_hd__conb_1 conb_T31Y47 (.HI(tie_high_T31Y47), .LO(tie_low_T31Y47));
  sky130_fd_sc_hd__conb_1 conb_T31Y48 (.HI(tie_high_T31Y48), .LO(tie_low_T31Y48));
  sky130_fd_sc_hd__conb_1 conb_T31Y49 (.HI(tie_high_T31Y49), .LO(tie_low_T31Y49));
  sky130_fd_sc_hd__conb_1 conb_T31Y5 (.HI(tie_high_T31Y5), .LO(tie_low_T31Y5));
  sky130_fd_sc_hd__conb_1 conb_T31Y50 (.HI(tie_high_T31Y50), .LO(tie_low_T31Y50));
  sky130_fd_sc_hd__conb_1 conb_T31Y51 (.HI(tie_high_T31Y51), .LO(tie_low_T31Y51));
  sky130_fd_sc_hd__conb_1 conb_T31Y52 (.HI(tie_high_T31Y52), .LO(tie_low_T31Y52));
  sky130_fd_sc_hd__conb_1 conb_T31Y53 (.HI(tie_high_T31Y53), .LO(tie_low_T31Y53));
  sky130_fd_sc_hd__conb_1 conb_T31Y54 (.HI(tie_high_T31Y54), .LO(tie_low_T31Y54));
  sky130_fd_sc_hd__conb_1 conb_T31Y55 (.HI(tie_high_T31Y55), .LO(tie_low_T31Y55));
  sky130_fd_sc_hd__conb_1 conb_T31Y56 (.HI(tie_high_T31Y56), .LO(tie_low_T31Y56));
  sky130_fd_sc_hd__conb_1 conb_T31Y57 (.HI(tie_high_T31Y57), .LO(tie_low_T31Y57));
  sky130_fd_sc_hd__conb_1 conb_T31Y58 (.HI(tie_high_T31Y58), .LO(tie_low_T31Y58));
  sky130_fd_sc_hd__conb_1 conb_T31Y59 (.HI(tie_high_T31Y59), .LO(tie_low_T31Y59));
  sky130_fd_sc_hd__conb_1 conb_T31Y6 (.HI(tie_high_T31Y6), .LO(tie_low_T31Y6));
  sky130_fd_sc_hd__conb_1 conb_T31Y60 (.HI(tie_high_T31Y60), .LO(tie_low_T31Y60));
  sky130_fd_sc_hd__conb_1 conb_T31Y61 (.HI(tie_high_T31Y61), .LO(tie_low_T31Y61));
  sky130_fd_sc_hd__conb_1 conb_T31Y62 (.HI(tie_high_T31Y62), .LO(tie_low_T31Y62));
  sky130_fd_sc_hd__conb_1 conb_T31Y63 (.HI(tie_high_T31Y63), .LO(tie_low_T31Y63));
  sky130_fd_sc_hd__conb_1 conb_T31Y64 (.HI(tie_high_T31Y64), .LO(tie_low_T31Y64));
  sky130_fd_sc_hd__conb_1 conb_T31Y65 (.HI(tie_high_T31Y65), .LO(tie_low_T31Y65));
  sky130_fd_sc_hd__conb_1 conb_T31Y66 (.HI(tie_high_T31Y66), .LO(tie_low_T31Y66));
  sky130_fd_sc_hd__conb_1 conb_T31Y67 (.HI(tie_high_T31Y67), .LO(tie_low_T31Y67));
  sky130_fd_sc_hd__conb_1 conb_T31Y68 (.HI(tie_high_T31Y68), .LO(tie_low_T31Y68));
  sky130_fd_sc_hd__conb_1 conb_T31Y69 (.HI(tie_high_T31Y69), .LO(tie_low_T31Y69));
  sky130_fd_sc_hd__conb_1 conb_T31Y7 (.HI(tie_high_T31Y7), .LO(tie_low_T31Y7));
  sky130_fd_sc_hd__conb_1 conb_T31Y70 (.HI(tie_high_T31Y70), .LO(tie_low_T31Y70));
  sky130_fd_sc_hd__conb_1 conb_T31Y71 (.HI(tie_high_T31Y71), .LO(tie_low_T31Y71));
  sky130_fd_sc_hd__conb_1 conb_T31Y72 (.HI(tie_high_T31Y72), .LO(tie_low_T31Y72));
  sky130_fd_sc_hd__conb_1 conb_T31Y73 (.HI(tie_high_T31Y73), .LO(tie_low_T31Y73));
  sky130_fd_sc_hd__conb_1 conb_T31Y74 (.HI(tie_high_T31Y74), .LO(tie_low_T31Y74));
  sky130_fd_sc_hd__conb_1 conb_T31Y75 (.HI(tie_high_T31Y75), .LO(tie_low_T31Y75));
  sky130_fd_sc_hd__conb_1 conb_T31Y76 (.HI(tie_high_T31Y76), .LO(tie_low_T31Y76));
  sky130_fd_sc_hd__conb_1 conb_T31Y77 (.HI(tie_high_T31Y77), .LO(tie_low_T31Y77));
  sky130_fd_sc_hd__conb_1 conb_T31Y78 (.HI(tie_high_T31Y78), .LO(tie_low_T31Y78));
  sky130_fd_sc_hd__conb_1 conb_T31Y79 (.HI(tie_high_T31Y79), .LO(tie_low_T31Y79));
  sky130_fd_sc_hd__conb_1 conb_T31Y8 (.HI(tie_high_T31Y8), .LO(tie_low_T31Y8));
  sky130_fd_sc_hd__conb_1 conb_T31Y80 (.HI(tie_high_T31Y80), .LO(tie_low_T31Y80));
  sky130_fd_sc_hd__conb_1 conb_T31Y81 (.HI(tie_high_T31Y81), .LO(tie_low_T31Y81));
  sky130_fd_sc_hd__conb_1 conb_T31Y82 (.HI(tie_high_T31Y82), .LO(tie_low_T31Y82));
  sky130_fd_sc_hd__conb_1 conb_T31Y83 (.HI(tie_high_T31Y83), .LO(tie_low_T31Y83));
  sky130_fd_sc_hd__conb_1 conb_T31Y84 (.HI(tie_high_T31Y84), .LO(tie_low_T31Y84));
  sky130_fd_sc_hd__conb_1 conb_T31Y85 (.HI(tie_high_T31Y85), .LO(tie_low_T31Y85));
  sky130_fd_sc_hd__conb_1 conb_T31Y86 (.HI(tie_high_T31Y86), .LO(tie_low_T31Y86));
  sky130_fd_sc_hd__conb_1 conb_T31Y87 (.HI(tie_high_T31Y87), .LO(tie_low_T31Y87));
  sky130_fd_sc_hd__conb_1 conb_T31Y88 (.HI(tie_high_T31Y88), .LO(tie_low_T31Y88));
  sky130_fd_sc_hd__conb_1 conb_T31Y89 (.HI(tie_high_T31Y89), .LO(tie_low_T31Y89));
  sky130_fd_sc_hd__conb_1 conb_T31Y9 (.HI(tie_high_T31Y9), .LO(tie_low_T31Y9));
  sky130_fd_sc_hd__conb_1 conb_T32Y0 (.HI(tie_high_T32Y0), .LO(tie_low_T32Y0));
  sky130_fd_sc_hd__conb_1 conb_T32Y1 (.HI(tie_high_T32Y1), .LO(tie_low_T32Y1));
  sky130_fd_sc_hd__conb_1 conb_T32Y10 (.HI(tie_high_T32Y10), .LO(tie_low_T32Y10));
  sky130_fd_sc_hd__conb_1 conb_T32Y11 (.HI(tie_high_T32Y11), .LO(tie_low_T32Y11));
  sky130_fd_sc_hd__conb_1 conb_T32Y12 (.HI(tie_high_T32Y12), .LO(tie_low_T32Y12));
  sky130_fd_sc_hd__conb_1 conb_T32Y13 (.HI(tie_high_T32Y13), .LO(tie_low_T32Y13));
  sky130_fd_sc_hd__conb_1 conb_T32Y14 (.HI(tie_high_T32Y14), .LO(tie_low_T32Y14));
  sky130_fd_sc_hd__conb_1 conb_T32Y15 (.HI(tie_high_T32Y15), .LO(tie_low_T32Y15));
  sky130_fd_sc_hd__conb_1 conb_T32Y16 (.HI(tie_high_T32Y16), .LO(tie_low_T32Y16));
  sky130_fd_sc_hd__conb_1 conb_T32Y17 (.HI(tie_high_T32Y17), .LO(tie_low_T32Y17));
  sky130_fd_sc_hd__conb_1 conb_T32Y18 (.HI(tie_high_T32Y18), .LO(tie_low_T32Y18));
  sky130_fd_sc_hd__conb_1 conb_T32Y19 (.HI(tie_high_T32Y19), .LO(tie_low_T32Y19));
  sky130_fd_sc_hd__conb_1 conb_T32Y2 (.HI(tie_high_T32Y2), .LO(tie_low_T32Y2));
  sky130_fd_sc_hd__conb_1 conb_T32Y20 (.HI(tie_high_T32Y20), .LO(tie_low_T32Y20));
  sky130_fd_sc_hd__conb_1 conb_T32Y21 (.HI(tie_high_T32Y21), .LO(tie_low_T32Y21));
  sky130_fd_sc_hd__conb_1 conb_T32Y22 (.HI(tie_high_T32Y22), .LO(tie_low_T32Y22));
  sky130_fd_sc_hd__conb_1 conb_T32Y23 (.HI(tie_high_T32Y23), .LO(tie_low_T32Y23));
  sky130_fd_sc_hd__conb_1 conb_T32Y24 (.HI(tie_high_T32Y24), .LO(tie_low_T32Y24));
  sky130_fd_sc_hd__conb_1 conb_T32Y25 (.HI(tie_high_T32Y25), .LO(tie_low_T32Y25));
  sky130_fd_sc_hd__conb_1 conb_T32Y26 (.HI(tie_high_T32Y26), .LO(tie_low_T32Y26));
  sky130_fd_sc_hd__conb_1 conb_T32Y27 (.HI(tie_high_T32Y27), .LO(tie_low_T32Y27));
  sky130_fd_sc_hd__conb_1 conb_T32Y28 (.HI(tie_high_T32Y28), .LO(tie_low_T32Y28));
  sky130_fd_sc_hd__conb_1 conb_T32Y29 (.HI(tie_high_T32Y29), .LO(tie_low_T32Y29));
  sky130_fd_sc_hd__conb_1 conb_T32Y3 (.HI(tie_high_T32Y3), .LO(tie_low_T32Y3));
  sky130_fd_sc_hd__conb_1 conb_T32Y30 (.HI(tie_high_T32Y30), .LO(tie_low_T32Y30));
  sky130_fd_sc_hd__conb_1 conb_T32Y31 (.HI(tie_high_T32Y31), .LO(tie_low_T32Y31));
  sky130_fd_sc_hd__conb_1 conb_T32Y32 (.HI(tie_high_T32Y32), .LO(tie_low_T32Y32));
  sky130_fd_sc_hd__conb_1 conb_T32Y33 (.HI(tie_high_T32Y33), .LO(tie_low_T32Y33));
  sky130_fd_sc_hd__conb_1 conb_T32Y34 (.HI(tie_high_T32Y34), .LO(tie_low_T32Y34));
  sky130_fd_sc_hd__conb_1 conb_T32Y35 (.HI(tie_high_T32Y35), .LO(tie_low_T32Y35));
  sky130_fd_sc_hd__conb_1 conb_T32Y36 (.HI(tie_high_T32Y36), .LO(tie_low_T32Y36));
  sky130_fd_sc_hd__conb_1 conb_T32Y37 (.HI(tie_high_T32Y37), .LO(tie_low_T32Y37));
  sky130_fd_sc_hd__conb_1 conb_T32Y38 (.HI(tie_high_T32Y38), .LO(tie_low_T32Y38));
  sky130_fd_sc_hd__conb_1 conb_T32Y39 (.HI(tie_high_T32Y39), .LO(tie_low_T32Y39));
  sky130_fd_sc_hd__conb_1 conb_T32Y4 (.HI(tie_high_T32Y4), .LO(tie_low_T32Y4));
  sky130_fd_sc_hd__conb_1 conb_T32Y40 (.HI(tie_high_T32Y40), .LO(tie_low_T32Y40));
  sky130_fd_sc_hd__conb_1 conb_T32Y41 (.HI(tie_high_T32Y41), .LO(tie_low_T32Y41));
  sky130_fd_sc_hd__conb_1 conb_T32Y42 (.HI(tie_high_T32Y42), .LO(tie_low_T32Y42));
  sky130_fd_sc_hd__conb_1 conb_T32Y43 (.HI(tie_high_T32Y43), .LO(tie_low_T32Y43));
  sky130_fd_sc_hd__conb_1 conb_T32Y44 (.HI(tie_high_T32Y44), .LO(tie_low_T32Y44));
  sky130_fd_sc_hd__conb_1 conb_T32Y45 (.HI(tie_high_T32Y45), .LO(tie_low_T32Y45));
  sky130_fd_sc_hd__conb_1 conb_T32Y46 (.HI(tie_high_T32Y46), .LO(tie_low_T32Y46));
  sky130_fd_sc_hd__conb_1 conb_T32Y47 (.HI(tie_high_T32Y47), .LO(tie_low_T32Y47));
  sky130_fd_sc_hd__conb_1 conb_T32Y48 (.HI(tie_high_T32Y48), .LO(tie_low_T32Y48));
  sky130_fd_sc_hd__conb_1 conb_T32Y49 (.HI(tie_high_T32Y49), .LO(tie_low_T32Y49));
  sky130_fd_sc_hd__conb_1 conb_T32Y5 (.HI(tie_high_T32Y5), .LO(tie_low_T32Y5));
  sky130_fd_sc_hd__conb_1 conb_T32Y50 (.HI(tie_high_T32Y50), .LO(tie_low_T32Y50));
  sky130_fd_sc_hd__conb_1 conb_T32Y51 (.HI(tie_high_T32Y51), .LO(tie_low_T32Y51));
  sky130_fd_sc_hd__conb_1 conb_T32Y52 (.HI(tie_high_T32Y52), .LO(tie_low_T32Y52));
  sky130_fd_sc_hd__conb_1 conb_T32Y53 (.HI(tie_high_T32Y53), .LO(tie_low_T32Y53));
  sky130_fd_sc_hd__conb_1 conb_T32Y54 (.HI(tie_high_T32Y54), .LO(tie_low_T32Y54));
  sky130_fd_sc_hd__conb_1 conb_T32Y55 (.HI(tie_high_T32Y55), .LO(tie_low_T32Y55));
  sky130_fd_sc_hd__conb_1 conb_T32Y56 (.HI(tie_high_T32Y56), .LO(tie_low_T32Y56));
  sky130_fd_sc_hd__conb_1 conb_T32Y57 (.HI(tie_high_T32Y57), .LO(tie_low_T32Y57));
  sky130_fd_sc_hd__conb_1 conb_T32Y58 (.HI(tie_high_T32Y58), .LO(tie_low_T32Y58));
  sky130_fd_sc_hd__conb_1 conb_T32Y59 (.HI(tie_high_T32Y59), .LO(tie_low_T32Y59));
  sky130_fd_sc_hd__conb_1 conb_T32Y6 (.HI(tie_high_T32Y6), .LO(tie_low_T32Y6));
  sky130_fd_sc_hd__conb_1 conb_T32Y60 (.HI(tie_high_T32Y60), .LO(tie_low_T32Y60));
  sky130_fd_sc_hd__conb_1 conb_T32Y61 (.HI(tie_high_T32Y61), .LO(tie_low_T32Y61));
  sky130_fd_sc_hd__conb_1 conb_T32Y62 (.HI(tie_high_T32Y62), .LO(tie_low_T32Y62));
  sky130_fd_sc_hd__conb_1 conb_T32Y63 (.HI(tie_high_T32Y63), .LO(tie_low_T32Y63));
  sky130_fd_sc_hd__conb_1 conb_T32Y64 (.HI(tie_high_T32Y64), .LO(tie_low_T32Y64));
  sky130_fd_sc_hd__conb_1 conb_T32Y65 (.HI(tie_high_T32Y65), .LO(tie_low_T32Y65));
  sky130_fd_sc_hd__conb_1 conb_T32Y66 (.HI(tie_high_T32Y66), .LO(tie_low_T32Y66));
  sky130_fd_sc_hd__conb_1 conb_T32Y67 (.HI(tie_high_T32Y67), .LO(tie_low_T32Y67));
  sky130_fd_sc_hd__conb_1 conb_T32Y68 (.HI(tie_high_T32Y68), .LO(tie_low_T32Y68));
  sky130_fd_sc_hd__conb_1 conb_T32Y69 (.HI(tie_high_T32Y69), .LO(tie_low_T32Y69));
  sky130_fd_sc_hd__conb_1 conb_T32Y7 (.HI(tie_high_T32Y7), .LO(tie_low_T32Y7));
  sky130_fd_sc_hd__conb_1 conb_T32Y70 (.HI(tie_high_T32Y70), .LO(tie_low_T32Y70));
  sky130_fd_sc_hd__conb_1 conb_T32Y71 (.HI(tie_high_T32Y71), .LO(tie_low_T32Y71));
  sky130_fd_sc_hd__conb_1 conb_T32Y72 (.HI(tie_high_T32Y72), .LO(tie_low_T32Y72));
  sky130_fd_sc_hd__conb_1 conb_T32Y73 (.HI(tie_high_T32Y73), .LO(tie_low_T32Y73));
  sky130_fd_sc_hd__conb_1 conb_T32Y74 (.HI(tie_high_T32Y74), .LO(tie_low_T32Y74));
  sky130_fd_sc_hd__conb_1 conb_T32Y75 (.HI(tie_high_T32Y75), .LO(tie_low_T32Y75));
  sky130_fd_sc_hd__conb_1 conb_T32Y76 (.HI(tie_high_T32Y76), .LO(tie_low_T32Y76));
  sky130_fd_sc_hd__conb_1 conb_T32Y77 (.HI(tie_high_T32Y77), .LO(tie_low_T32Y77));
  sky130_fd_sc_hd__conb_1 conb_T32Y78 (.HI(tie_high_T32Y78), .LO(tie_low_T32Y78));
  sky130_fd_sc_hd__conb_1 conb_T32Y79 (.HI(tie_high_T32Y79), .LO(tie_low_T32Y79));
  sky130_fd_sc_hd__conb_1 conb_T32Y8 (.HI(tie_high_T32Y8), .LO(tie_low_T32Y8));
  sky130_fd_sc_hd__conb_1 conb_T32Y80 (.HI(tie_high_T32Y80), .LO(tie_low_T32Y80));
  sky130_fd_sc_hd__conb_1 conb_T32Y81 (.HI(tie_high_T32Y81), .LO(tie_low_T32Y81));
  sky130_fd_sc_hd__conb_1 conb_T32Y82 (.HI(tie_high_T32Y82), .LO(tie_low_T32Y82));
  sky130_fd_sc_hd__conb_1 conb_T32Y83 (.HI(tie_high_T32Y83), .LO(tie_low_T32Y83));
  sky130_fd_sc_hd__conb_1 conb_T32Y84 (.HI(tie_high_T32Y84), .LO(tie_low_T32Y84));
  sky130_fd_sc_hd__conb_1 conb_T32Y85 (.HI(tie_high_T32Y85), .LO(tie_low_T32Y85));
  sky130_fd_sc_hd__conb_1 conb_T32Y86 (.HI(tie_high_T32Y86), .LO(tie_low_T32Y86));
  sky130_fd_sc_hd__conb_1 conb_T32Y87 (.HI(tie_high_T32Y87), .LO(tie_low_T32Y87));
  sky130_fd_sc_hd__conb_1 conb_T32Y88 (.HI(tie_high_T32Y88), .LO(tie_low_T32Y88));
  sky130_fd_sc_hd__conb_1 conb_T32Y89 (.HI(tie_high_T32Y89), .LO(tie_low_T32Y89));
  sky130_fd_sc_hd__conb_1 conb_T32Y9 (.HI(tie_high_T32Y9), .LO(tie_low_T32Y9));
  sky130_fd_sc_hd__conb_1 conb_T33Y0 (.HI(tie_high_T33Y0), .LO(tie_low_T33Y0));
  sky130_fd_sc_hd__conb_1 conb_T33Y1 (.HI(tie_high_T33Y1), .LO(tie_low_T33Y1));
  sky130_fd_sc_hd__conb_1 conb_T33Y10 (.HI(tie_high_T33Y10), .LO(tie_low_T33Y10));
  sky130_fd_sc_hd__conb_1 conb_T33Y11 (.HI(tie_high_T33Y11), .LO(tie_low_T33Y11));
  sky130_fd_sc_hd__conb_1 conb_T33Y12 (.HI(tie_high_T33Y12), .LO(tie_low_T33Y12));
  sky130_fd_sc_hd__conb_1 conb_T33Y13 (.HI(tie_high_T33Y13), .LO(tie_low_T33Y13));
  sky130_fd_sc_hd__conb_1 conb_T33Y14 (.HI(tie_high_T33Y14), .LO(tie_low_T33Y14));
  sky130_fd_sc_hd__conb_1 conb_T33Y15 (.HI(tie_high_T33Y15), .LO(tie_low_T33Y15));
  sky130_fd_sc_hd__conb_1 conb_T33Y16 (.HI(tie_high_T33Y16), .LO(tie_low_T33Y16));
  sky130_fd_sc_hd__conb_1 conb_T33Y17 (.HI(tie_high_T33Y17), .LO(tie_low_T33Y17));
  sky130_fd_sc_hd__conb_1 conb_T33Y18 (.HI(tie_high_T33Y18), .LO(tie_low_T33Y18));
  sky130_fd_sc_hd__conb_1 conb_T33Y19 (.HI(tie_high_T33Y19), .LO(tie_low_T33Y19));
  sky130_fd_sc_hd__conb_1 conb_T33Y2 (.HI(tie_high_T33Y2), .LO(tie_low_T33Y2));
  sky130_fd_sc_hd__conb_1 conb_T33Y20 (.HI(tie_high_T33Y20), .LO(tie_low_T33Y20));
  sky130_fd_sc_hd__conb_1 conb_T33Y21 (.HI(tie_high_T33Y21), .LO(tie_low_T33Y21));
  sky130_fd_sc_hd__conb_1 conb_T33Y22 (.HI(tie_high_T33Y22), .LO(tie_low_T33Y22));
  sky130_fd_sc_hd__conb_1 conb_T33Y23 (.HI(tie_high_T33Y23), .LO(tie_low_T33Y23));
  sky130_fd_sc_hd__conb_1 conb_T33Y24 (.HI(tie_high_T33Y24), .LO(tie_low_T33Y24));
  sky130_fd_sc_hd__conb_1 conb_T33Y25 (.HI(tie_high_T33Y25), .LO(tie_low_T33Y25));
  sky130_fd_sc_hd__conb_1 conb_T33Y26 (.HI(tie_high_T33Y26), .LO(tie_low_T33Y26));
  sky130_fd_sc_hd__conb_1 conb_T33Y27 (.HI(tie_high_T33Y27), .LO(tie_low_T33Y27));
  sky130_fd_sc_hd__conb_1 conb_T33Y28 (.HI(tie_high_T33Y28), .LO(tie_low_T33Y28));
  sky130_fd_sc_hd__conb_1 conb_T33Y29 (.HI(tie_high_T33Y29), .LO(tie_low_T33Y29));
  sky130_fd_sc_hd__conb_1 conb_T33Y3 (.HI(tie_high_T33Y3), .LO(tie_low_T33Y3));
  sky130_fd_sc_hd__conb_1 conb_T33Y30 (.HI(tie_high_T33Y30), .LO(tie_low_T33Y30));
  sky130_fd_sc_hd__conb_1 conb_T33Y31 (.HI(tie_high_T33Y31), .LO(tie_low_T33Y31));
  sky130_fd_sc_hd__conb_1 conb_T33Y32 (.HI(tie_high_T33Y32), .LO(tie_low_T33Y32));
  sky130_fd_sc_hd__conb_1 conb_T33Y33 (.HI(tie_high_T33Y33), .LO(tie_low_T33Y33));
  sky130_fd_sc_hd__conb_1 conb_T33Y34 (.HI(tie_high_T33Y34), .LO(tie_low_T33Y34));
  sky130_fd_sc_hd__conb_1 conb_T33Y35 (.HI(tie_high_T33Y35), .LO(tie_low_T33Y35));
  sky130_fd_sc_hd__conb_1 conb_T33Y36 (.HI(tie_high_T33Y36), .LO(tie_low_T33Y36));
  sky130_fd_sc_hd__conb_1 conb_T33Y37 (.HI(tie_high_T33Y37), .LO(tie_low_T33Y37));
  sky130_fd_sc_hd__conb_1 conb_T33Y38 (.HI(tie_high_T33Y38), .LO(tie_low_T33Y38));
  sky130_fd_sc_hd__conb_1 conb_T33Y39 (.HI(tie_high_T33Y39), .LO(tie_low_T33Y39));
  sky130_fd_sc_hd__conb_1 conb_T33Y4 (.HI(tie_high_T33Y4), .LO(tie_low_T33Y4));
  sky130_fd_sc_hd__conb_1 conb_T33Y40 (.HI(tie_high_T33Y40), .LO(tie_low_T33Y40));
  sky130_fd_sc_hd__conb_1 conb_T33Y41 (.HI(tie_high_T33Y41), .LO(tie_low_T33Y41));
  sky130_fd_sc_hd__conb_1 conb_T33Y42 (.HI(tie_high_T33Y42), .LO(tie_low_T33Y42));
  sky130_fd_sc_hd__conb_1 conb_T33Y43 (.HI(tie_high_T33Y43), .LO(tie_low_T33Y43));
  sky130_fd_sc_hd__conb_1 conb_T33Y44 (.HI(tie_high_T33Y44), .LO(tie_low_T33Y44));
  sky130_fd_sc_hd__conb_1 conb_T33Y45 (.HI(tie_high_T33Y45), .LO(tie_low_T33Y45));
  sky130_fd_sc_hd__conb_1 conb_T33Y46 (.HI(tie_high_T33Y46), .LO(tie_low_T33Y46));
  sky130_fd_sc_hd__conb_1 conb_T33Y47 (.HI(tie_high_T33Y47), .LO(tie_low_T33Y47));
  sky130_fd_sc_hd__conb_1 conb_T33Y48 (.HI(tie_high_T33Y48), .LO(tie_low_T33Y48));
  sky130_fd_sc_hd__conb_1 conb_T33Y49 (.HI(tie_high_T33Y49), .LO(tie_low_T33Y49));
  sky130_fd_sc_hd__conb_1 conb_T33Y5 (.HI(tie_high_T33Y5), .LO(tie_low_T33Y5));
  sky130_fd_sc_hd__conb_1 conb_T33Y50 (.HI(tie_high_T33Y50), .LO(tie_low_T33Y50));
  sky130_fd_sc_hd__conb_1 conb_T33Y51 (.HI(tie_high_T33Y51), .LO(tie_low_T33Y51));
  sky130_fd_sc_hd__conb_1 conb_T33Y52 (.HI(tie_high_T33Y52), .LO(tie_low_T33Y52));
  sky130_fd_sc_hd__conb_1 conb_T33Y53 (.HI(tie_high_T33Y53), .LO(tie_low_T33Y53));
  sky130_fd_sc_hd__conb_1 conb_T33Y54 (.HI(tie_high_T33Y54), .LO(tie_low_T33Y54));
  sky130_fd_sc_hd__conb_1 conb_T33Y55 (.HI(tie_high_T33Y55), .LO(tie_low_T33Y55));
  sky130_fd_sc_hd__conb_1 conb_T33Y56 (.HI(tie_high_T33Y56), .LO(tie_low_T33Y56));
  sky130_fd_sc_hd__conb_1 conb_T33Y57 (.HI(tie_high_T33Y57), .LO(tie_low_T33Y57));
  sky130_fd_sc_hd__conb_1 conb_T33Y58 (.HI(tie_high_T33Y58), .LO(tie_low_T33Y58));
  sky130_fd_sc_hd__conb_1 conb_T33Y59 (.HI(tie_high_T33Y59), .LO(tie_low_T33Y59));
  sky130_fd_sc_hd__conb_1 conb_T33Y6 (.HI(tie_high_T33Y6), .LO(tie_low_T33Y6));
  sky130_fd_sc_hd__conb_1 conb_T33Y60 (.HI(tie_high_T33Y60), .LO(tie_low_T33Y60));
  sky130_fd_sc_hd__conb_1 conb_T33Y61 (.HI(tie_high_T33Y61), .LO(tie_low_T33Y61));
  sky130_fd_sc_hd__conb_1 conb_T33Y62 (.HI(tie_high_T33Y62), .LO(tie_low_T33Y62));
  sky130_fd_sc_hd__conb_1 conb_T33Y63 (.HI(tie_high_T33Y63), .LO(tie_low_T33Y63));
  sky130_fd_sc_hd__conb_1 conb_T33Y64 (.HI(tie_high_T33Y64), .LO(tie_low_T33Y64));
  sky130_fd_sc_hd__conb_1 conb_T33Y65 (.HI(tie_high_T33Y65), .LO(tie_low_T33Y65));
  sky130_fd_sc_hd__conb_1 conb_T33Y66 (.HI(tie_high_T33Y66), .LO(tie_low_T33Y66));
  sky130_fd_sc_hd__conb_1 conb_T33Y67 (.HI(tie_high_T33Y67), .LO(tie_low_T33Y67));
  sky130_fd_sc_hd__conb_1 conb_T33Y68 (.HI(tie_high_T33Y68), .LO(tie_low_T33Y68));
  sky130_fd_sc_hd__conb_1 conb_T33Y69 (.HI(tie_high_T33Y69), .LO(tie_low_T33Y69));
  sky130_fd_sc_hd__conb_1 conb_T33Y7 (.HI(tie_high_T33Y7), .LO(tie_low_T33Y7));
  sky130_fd_sc_hd__conb_1 conb_T33Y70 (.HI(tie_high_T33Y70), .LO(tie_low_T33Y70));
  sky130_fd_sc_hd__conb_1 conb_T33Y71 (.HI(tie_high_T33Y71), .LO(tie_low_T33Y71));
  sky130_fd_sc_hd__conb_1 conb_T33Y72 (.HI(tie_high_T33Y72), .LO(tie_low_T33Y72));
  sky130_fd_sc_hd__conb_1 conb_T33Y73 (.HI(tie_high_T33Y73), .LO(tie_low_T33Y73));
  sky130_fd_sc_hd__conb_1 conb_T33Y74 (.HI(tie_high_T33Y74), .LO(tie_low_T33Y74));
  sky130_fd_sc_hd__conb_1 conb_T33Y75 (.HI(tie_high_T33Y75), .LO(tie_low_T33Y75));
  sky130_fd_sc_hd__conb_1 conb_T33Y76 (.HI(tie_high_T33Y76), .LO(tie_low_T33Y76));
  sky130_fd_sc_hd__conb_1 conb_T33Y77 (.HI(tie_high_T33Y77), .LO(tie_low_T33Y77));
  sky130_fd_sc_hd__conb_1 conb_T33Y78 (.HI(tie_high_T33Y78), .LO(tie_low_T33Y78));
  sky130_fd_sc_hd__conb_1 conb_T33Y79 (.HI(tie_high_T33Y79), .LO(tie_low_T33Y79));
  sky130_fd_sc_hd__conb_1 conb_T33Y8 (.HI(tie_high_T33Y8), .LO(tie_low_T33Y8));
  sky130_fd_sc_hd__conb_1 conb_T33Y80 (.HI(tie_high_T33Y80), .LO(tie_low_T33Y80));
  sky130_fd_sc_hd__conb_1 conb_T33Y81 (.HI(tie_high_T33Y81), .LO(tie_low_T33Y81));
  sky130_fd_sc_hd__conb_1 conb_T33Y82 (.HI(tie_high_T33Y82), .LO(tie_low_T33Y82));
  sky130_fd_sc_hd__conb_1 conb_T33Y83 (.HI(tie_high_T33Y83), .LO(tie_low_T33Y83));
  sky130_fd_sc_hd__conb_1 conb_T33Y84 (.HI(tie_high_T33Y84), .LO(tie_low_T33Y84));
  sky130_fd_sc_hd__conb_1 conb_T33Y85 (.HI(tie_high_T33Y85), .LO(tie_low_T33Y85));
  sky130_fd_sc_hd__conb_1 conb_T33Y86 (.HI(tie_high_T33Y86), .LO(tie_low_T33Y86));
  sky130_fd_sc_hd__conb_1 conb_T33Y87 (.HI(tie_high_T33Y87), .LO(tie_low_T33Y87));
  sky130_fd_sc_hd__conb_1 conb_T33Y88 (.HI(tie_high_T33Y88), .LO(tie_low_T33Y88));
  sky130_fd_sc_hd__conb_1 conb_T33Y89 (.HI(tie_high_T33Y89), .LO(tie_low_T33Y89));
  sky130_fd_sc_hd__conb_1 conb_T33Y9 (.HI(tie_high_T33Y9), .LO(tie_low_T33Y9));
  sky130_fd_sc_hd__conb_1 conb_T34Y0 (.HI(tie_high_T34Y0), .LO(tie_low_T34Y0));
  sky130_fd_sc_hd__conb_1 conb_T34Y1 (.HI(tie_high_T34Y1), .LO(tie_low_T34Y1));
  sky130_fd_sc_hd__conb_1 conb_T34Y10 (.HI(tie_high_T34Y10), .LO(tie_low_T34Y10));
  sky130_fd_sc_hd__conb_1 conb_T34Y11 (.HI(tie_high_T34Y11), .LO(tie_low_T34Y11));
  sky130_fd_sc_hd__conb_1 conb_T34Y12 (.HI(tie_high_T34Y12), .LO(tie_low_T34Y12));
  sky130_fd_sc_hd__conb_1 conb_T34Y13 (.HI(tie_high_T34Y13), .LO(tie_low_T34Y13));
  sky130_fd_sc_hd__conb_1 conb_T34Y14 (.HI(tie_high_T34Y14), .LO(tie_low_T34Y14));
  sky130_fd_sc_hd__conb_1 conb_T34Y15 (.HI(tie_high_T34Y15), .LO(tie_low_T34Y15));
  sky130_fd_sc_hd__conb_1 conb_T34Y16 (.HI(tie_high_T34Y16), .LO(tie_low_T34Y16));
  sky130_fd_sc_hd__conb_1 conb_T34Y17 (.HI(tie_high_T34Y17), .LO(tie_low_T34Y17));
  sky130_fd_sc_hd__conb_1 conb_T34Y18 (.HI(tie_high_T34Y18), .LO(tie_low_T34Y18));
  sky130_fd_sc_hd__conb_1 conb_T34Y19 (.HI(tie_high_T34Y19), .LO(tie_low_T34Y19));
  sky130_fd_sc_hd__conb_1 conb_T34Y2 (.HI(tie_high_T34Y2), .LO(tie_low_T34Y2));
  sky130_fd_sc_hd__conb_1 conb_T34Y20 (.HI(tie_high_T34Y20), .LO(tie_low_T34Y20));
  sky130_fd_sc_hd__conb_1 conb_T34Y21 (.HI(tie_high_T34Y21), .LO(tie_low_T34Y21));
  sky130_fd_sc_hd__conb_1 conb_T34Y22 (.HI(tie_high_T34Y22), .LO(tie_low_T34Y22));
  sky130_fd_sc_hd__conb_1 conb_T34Y23 (.HI(tie_high_T34Y23), .LO(tie_low_T34Y23));
  sky130_fd_sc_hd__conb_1 conb_T34Y24 (.HI(tie_high_T34Y24), .LO(tie_low_T34Y24));
  sky130_fd_sc_hd__conb_1 conb_T34Y25 (.HI(tie_high_T34Y25), .LO(tie_low_T34Y25));
  sky130_fd_sc_hd__conb_1 conb_T34Y26 (.HI(tie_high_T34Y26), .LO(tie_low_T34Y26));
  sky130_fd_sc_hd__conb_1 conb_T34Y27 (.HI(tie_high_T34Y27), .LO(tie_low_T34Y27));
  sky130_fd_sc_hd__conb_1 conb_T34Y28 (.HI(tie_high_T34Y28), .LO(tie_low_T34Y28));
  sky130_fd_sc_hd__conb_1 conb_T34Y29 (.HI(tie_high_T34Y29), .LO(tie_low_T34Y29));
  sky130_fd_sc_hd__conb_1 conb_T34Y3 (.HI(tie_high_T34Y3), .LO(tie_low_T34Y3));
  sky130_fd_sc_hd__conb_1 conb_T34Y30 (.HI(tie_high_T34Y30), .LO(tie_low_T34Y30));
  sky130_fd_sc_hd__conb_1 conb_T34Y31 (.HI(tie_high_T34Y31), .LO(tie_low_T34Y31));
  sky130_fd_sc_hd__conb_1 conb_T34Y32 (.HI(tie_high_T34Y32), .LO(tie_low_T34Y32));
  sky130_fd_sc_hd__conb_1 conb_T34Y33 (.HI(tie_high_T34Y33), .LO(tie_low_T34Y33));
  sky130_fd_sc_hd__conb_1 conb_T34Y34 (.HI(tie_high_T34Y34), .LO(tie_low_T34Y34));
  sky130_fd_sc_hd__conb_1 conb_T34Y35 (.HI(tie_high_T34Y35), .LO(tie_low_T34Y35));
  sky130_fd_sc_hd__conb_1 conb_T34Y36 (.HI(tie_high_T34Y36), .LO(tie_low_T34Y36));
  sky130_fd_sc_hd__conb_1 conb_T34Y37 (.HI(tie_high_T34Y37), .LO(tie_low_T34Y37));
  sky130_fd_sc_hd__conb_1 conb_T34Y38 (.HI(tie_high_T34Y38), .LO(tie_low_T34Y38));
  sky130_fd_sc_hd__conb_1 conb_T34Y39 (.HI(tie_high_T34Y39), .LO(tie_low_T34Y39));
  sky130_fd_sc_hd__conb_1 conb_T34Y4 (.HI(tie_high_T34Y4), .LO(tie_low_T34Y4));
  sky130_fd_sc_hd__conb_1 conb_T34Y40 (.HI(tie_high_T34Y40), .LO(tie_low_T34Y40));
  sky130_fd_sc_hd__conb_1 conb_T34Y41 (.HI(tie_high_T34Y41), .LO(tie_low_T34Y41));
  sky130_fd_sc_hd__conb_1 conb_T34Y42 (.HI(tie_high_T34Y42), .LO(tie_low_T34Y42));
  sky130_fd_sc_hd__conb_1 conb_T34Y43 (.HI(tie_high_T34Y43), .LO(tie_low_T34Y43));
  sky130_fd_sc_hd__conb_1 conb_T34Y44 (.HI(tie_high_T34Y44), .LO(tie_low_T34Y44));
  sky130_fd_sc_hd__conb_1 conb_T34Y45 (.HI(tie_high_T34Y45), .LO(tie_low_T34Y45));
  sky130_fd_sc_hd__conb_1 conb_T34Y46 (.HI(tie_high_T34Y46), .LO(tie_low_T34Y46));
  sky130_fd_sc_hd__conb_1 conb_T34Y47 (.HI(tie_high_T34Y47), .LO(tie_low_T34Y47));
  sky130_fd_sc_hd__conb_1 conb_T34Y48 (.HI(tie_high_T34Y48), .LO(tie_low_T34Y48));
  sky130_fd_sc_hd__conb_1 conb_T34Y49 (.HI(tie_high_T34Y49), .LO(tie_low_T34Y49));
  sky130_fd_sc_hd__conb_1 conb_T34Y5 (.HI(tie_high_T34Y5), .LO(tie_low_T34Y5));
  sky130_fd_sc_hd__conb_1 conb_T34Y50 (.HI(tie_high_T34Y50), .LO(tie_low_T34Y50));
  sky130_fd_sc_hd__conb_1 conb_T34Y51 (.HI(tie_high_T34Y51), .LO(tie_low_T34Y51));
  sky130_fd_sc_hd__conb_1 conb_T34Y52 (.HI(tie_high_T34Y52), .LO(tie_low_T34Y52));
  sky130_fd_sc_hd__conb_1 conb_T34Y53 (.HI(tie_high_T34Y53), .LO(tie_low_T34Y53));
  sky130_fd_sc_hd__conb_1 conb_T34Y54 (.HI(tie_high_T34Y54), .LO(tie_low_T34Y54));
  sky130_fd_sc_hd__conb_1 conb_T34Y55 (.HI(tie_high_T34Y55), .LO(tie_low_T34Y55));
  sky130_fd_sc_hd__conb_1 conb_T34Y56 (.HI(tie_high_T34Y56), .LO(tie_low_T34Y56));
  sky130_fd_sc_hd__conb_1 conb_T34Y57 (.HI(tie_high_T34Y57), .LO(tie_low_T34Y57));
  sky130_fd_sc_hd__conb_1 conb_T34Y58 (.HI(tie_high_T34Y58), .LO(tie_low_T34Y58));
  sky130_fd_sc_hd__conb_1 conb_T34Y59 (.HI(tie_high_T34Y59), .LO(tie_low_T34Y59));
  sky130_fd_sc_hd__conb_1 conb_T34Y6 (.HI(tie_high_T34Y6), .LO(tie_low_T34Y6));
  sky130_fd_sc_hd__conb_1 conb_T34Y60 (.HI(tie_high_T34Y60), .LO(tie_low_T34Y60));
  sky130_fd_sc_hd__conb_1 conb_T34Y61 (.HI(tie_high_T34Y61), .LO(tie_low_T34Y61));
  sky130_fd_sc_hd__conb_1 conb_T34Y62 (.HI(tie_high_T34Y62), .LO(tie_low_T34Y62));
  sky130_fd_sc_hd__conb_1 conb_T34Y63 (.HI(tie_high_T34Y63), .LO(tie_low_T34Y63));
  sky130_fd_sc_hd__conb_1 conb_T34Y64 (.HI(tie_high_T34Y64), .LO(tie_low_T34Y64));
  sky130_fd_sc_hd__conb_1 conb_T34Y65 (.HI(tie_high_T34Y65), .LO(tie_low_T34Y65));
  sky130_fd_sc_hd__conb_1 conb_T34Y66 (.HI(tie_high_T34Y66), .LO(tie_low_T34Y66));
  sky130_fd_sc_hd__conb_1 conb_T34Y67 (.HI(tie_high_T34Y67), .LO(tie_low_T34Y67));
  sky130_fd_sc_hd__conb_1 conb_T34Y68 (.HI(tie_high_T34Y68), .LO(tie_low_T34Y68));
  sky130_fd_sc_hd__conb_1 conb_T34Y69 (.HI(tie_high_T34Y69), .LO(tie_low_T34Y69));
  sky130_fd_sc_hd__conb_1 conb_T34Y7 (.HI(tie_high_T34Y7), .LO(tie_low_T34Y7));
  sky130_fd_sc_hd__conb_1 conb_T34Y70 (.HI(tie_high_T34Y70), .LO(tie_low_T34Y70));
  sky130_fd_sc_hd__conb_1 conb_T34Y71 (.HI(tie_high_T34Y71), .LO(tie_low_T34Y71));
  sky130_fd_sc_hd__conb_1 conb_T34Y72 (.HI(tie_high_T34Y72), .LO(tie_low_T34Y72));
  sky130_fd_sc_hd__conb_1 conb_T34Y73 (.HI(tie_high_T34Y73), .LO(tie_low_T34Y73));
  sky130_fd_sc_hd__conb_1 conb_T34Y74 (.HI(tie_high_T34Y74), .LO(tie_low_T34Y74));
  sky130_fd_sc_hd__conb_1 conb_T34Y75 (.HI(tie_high_T34Y75), .LO(tie_low_T34Y75));
  sky130_fd_sc_hd__conb_1 conb_T34Y76 (.HI(tie_high_T34Y76), .LO(tie_low_T34Y76));
  sky130_fd_sc_hd__conb_1 conb_T34Y77 (.HI(tie_high_T34Y77), .LO(tie_low_T34Y77));
  sky130_fd_sc_hd__conb_1 conb_T34Y78 (.HI(tie_high_T34Y78), .LO(tie_low_T34Y78));
  sky130_fd_sc_hd__conb_1 conb_T34Y79 (.HI(tie_high_T34Y79), .LO(tie_low_T34Y79));
  sky130_fd_sc_hd__conb_1 conb_T34Y8 (.HI(tie_high_T34Y8), .LO(tie_low_T34Y8));
  sky130_fd_sc_hd__conb_1 conb_T34Y80 (.HI(tie_high_T34Y80), .LO(tie_low_T34Y80));
  sky130_fd_sc_hd__conb_1 conb_T34Y81 (.HI(tie_high_T34Y81), .LO(tie_low_T34Y81));
  sky130_fd_sc_hd__conb_1 conb_T34Y82 (.HI(tie_high_T34Y82), .LO(tie_low_T34Y82));
  sky130_fd_sc_hd__conb_1 conb_T34Y83 (.HI(tie_high_T34Y83), .LO(tie_low_T34Y83));
  sky130_fd_sc_hd__conb_1 conb_T34Y84 (.HI(tie_high_T34Y84), .LO(tie_low_T34Y84));
  sky130_fd_sc_hd__conb_1 conb_T34Y85 (.HI(tie_high_T34Y85), .LO(tie_low_T34Y85));
  sky130_fd_sc_hd__conb_1 conb_T34Y86 (.HI(tie_high_T34Y86), .LO(tie_low_T34Y86));
  sky130_fd_sc_hd__conb_1 conb_T34Y87 (.HI(tie_high_T34Y87), .LO(tie_low_T34Y87));
  sky130_fd_sc_hd__conb_1 conb_T34Y88 (.HI(tie_high_T34Y88), .LO(tie_low_T34Y88));
  sky130_fd_sc_hd__conb_1 conb_T34Y89 (.HI(tie_high_T34Y89), .LO(tie_low_T34Y89));
  sky130_fd_sc_hd__conb_1 conb_T34Y9 (.HI(tie_high_T34Y9), .LO(tie_low_T34Y9));
  sky130_fd_sc_hd__conb_1 conb_T35Y0 (.HI(tie_high_T35Y0), .LO(tie_low_T35Y0));
  sky130_fd_sc_hd__conb_1 conb_T35Y1 (.HI(tie_high_T35Y1), .LO(tie_low_T35Y1));
  sky130_fd_sc_hd__conb_1 conb_T35Y10 (.HI(tie_high_T35Y10), .LO(tie_low_T35Y10));
  sky130_fd_sc_hd__conb_1 conb_T35Y11 (.HI(tie_high_T35Y11), .LO(tie_low_T35Y11));
  sky130_fd_sc_hd__conb_1 conb_T35Y12 (.HI(tie_high_T35Y12), .LO(tie_low_T35Y12));
  sky130_fd_sc_hd__conb_1 conb_T35Y13 (.HI(tie_high_T35Y13), .LO(tie_low_T35Y13));
  sky130_fd_sc_hd__conb_1 conb_T35Y14 (.HI(tie_high_T35Y14), .LO(tie_low_T35Y14));
  sky130_fd_sc_hd__conb_1 conb_T35Y15 (.HI(tie_high_T35Y15), .LO(tie_low_T35Y15));
  sky130_fd_sc_hd__conb_1 conb_T35Y16 (.HI(tie_high_T35Y16), .LO(tie_low_T35Y16));
  sky130_fd_sc_hd__conb_1 conb_T35Y17 (.HI(tie_high_T35Y17), .LO(tie_low_T35Y17));
  sky130_fd_sc_hd__conb_1 conb_T35Y18 (.HI(tie_high_T35Y18), .LO(tie_low_T35Y18));
  sky130_fd_sc_hd__conb_1 conb_T35Y19 (.HI(tie_high_T35Y19), .LO(tie_low_T35Y19));
  sky130_fd_sc_hd__conb_1 conb_T35Y2 (.HI(tie_high_T35Y2), .LO(tie_low_T35Y2));
  sky130_fd_sc_hd__conb_1 conb_T35Y20 (.HI(tie_high_T35Y20), .LO(tie_low_T35Y20));
  sky130_fd_sc_hd__conb_1 conb_T35Y21 (.HI(tie_high_T35Y21), .LO(tie_low_T35Y21));
  sky130_fd_sc_hd__conb_1 conb_T35Y22 (.HI(tie_high_T35Y22), .LO(tie_low_T35Y22));
  sky130_fd_sc_hd__conb_1 conb_T35Y23 (.HI(tie_high_T35Y23), .LO(tie_low_T35Y23));
  sky130_fd_sc_hd__conb_1 conb_T35Y24 (.HI(tie_high_T35Y24), .LO(tie_low_T35Y24));
  sky130_fd_sc_hd__conb_1 conb_T35Y25 (.HI(tie_high_T35Y25), .LO(tie_low_T35Y25));
  sky130_fd_sc_hd__conb_1 conb_T35Y26 (.HI(tie_high_T35Y26), .LO(tie_low_T35Y26));
  sky130_fd_sc_hd__conb_1 conb_T35Y27 (.HI(tie_high_T35Y27), .LO(tie_low_T35Y27));
  sky130_fd_sc_hd__conb_1 conb_T35Y28 (.HI(tie_high_T35Y28), .LO(tie_low_T35Y28));
  sky130_fd_sc_hd__conb_1 conb_T35Y29 (.HI(tie_high_T35Y29), .LO(tie_low_T35Y29));
  sky130_fd_sc_hd__conb_1 conb_T35Y3 (.HI(tie_high_T35Y3), .LO(tie_low_T35Y3));
  sky130_fd_sc_hd__conb_1 conb_T35Y30 (.HI(tie_high_T35Y30), .LO(tie_low_T35Y30));
  sky130_fd_sc_hd__conb_1 conb_T35Y31 (.HI(tie_high_T35Y31), .LO(tie_low_T35Y31));
  sky130_fd_sc_hd__conb_1 conb_T35Y32 (.HI(tie_high_T35Y32), .LO(tie_low_T35Y32));
  sky130_fd_sc_hd__conb_1 conb_T35Y33 (.HI(tie_high_T35Y33), .LO(tie_low_T35Y33));
  sky130_fd_sc_hd__conb_1 conb_T35Y34 (.HI(tie_high_T35Y34), .LO(tie_low_T35Y34));
  sky130_fd_sc_hd__conb_1 conb_T35Y35 (.HI(tie_high_T35Y35), .LO(tie_low_T35Y35));
  sky130_fd_sc_hd__conb_1 conb_T35Y36 (.HI(tie_high_T35Y36), .LO(tie_low_T35Y36));
  sky130_fd_sc_hd__conb_1 conb_T35Y37 (.HI(tie_high_T35Y37), .LO(tie_low_T35Y37));
  sky130_fd_sc_hd__conb_1 conb_T35Y38 (.HI(tie_high_T35Y38), .LO(tie_low_T35Y38));
  sky130_fd_sc_hd__conb_1 conb_T35Y39 (.HI(tie_high_T35Y39), .LO(tie_low_T35Y39));
  sky130_fd_sc_hd__conb_1 conb_T35Y4 (.HI(tie_high_T35Y4), .LO(tie_low_T35Y4));
  sky130_fd_sc_hd__conb_1 conb_T35Y40 (.HI(tie_high_T35Y40), .LO(tie_low_T35Y40));
  sky130_fd_sc_hd__conb_1 conb_T35Y41 (.HI(tie_high_T35Y41), .LO(tie_low_T35Y41));
  sky130_fd_sc_hd__conb_1 conb_T35Y42 (.HI(tie_high_T35Y42), .LO(tie_low_T35Y42));
  sky130_fd_sc_hd__conb_1 conb_T35Y43 (.HI(tie_high_T35Y43), .LO(tie_low_T35Y43));
  sky130_fd_sc_hd__conb_1 conb_T35Y44 (.HI(tie_high_T35Y44), .LO(tie_low_T35Y44));
  sky130_fd_sc_hd__conb_1 conb_T35Y45 (.HI(tie_high_T35Y45), .LO(tie_low_T35Y45));
  sky130_fd_sc_hd__conb_1 conb_T35Y46 (.HI(tie_high_T35Y46), .LO(tie_low_T35Y46));
  sky130_fd_sc_hd__conb_1 conb_T35Y47 (.HI(tie_high_T35Y47), .LO(tie_low_T35Y47));
  sky130_fd_sc_hd__conb_1 conb_T35Y48 (.HI(tie_high_T35Y48), .LO(tie_low_T35Y48));
  sky130_fd_sc_hd__conb_1 conb_T35Y49 (.HI(tie_high_T35Y49), .LO(tie_low_T35Y49));
  sky130_fd_sc_hd__conb_1 conb_T35Y5 (.HI(tie_high_T35Y5), .LO(tie_low_T35Y5));
  sky130_fd_sc_hd__conb_1 conb_T35Y50 (.HI(tie_high_T35Y50), .LO(tie_low_T35Y50));
  sky130_fd_sc_hd__conb_1 conb_T35Y51 (.HI(tie_high_T35Y51), .LO(tie_low_T35Y51));
  sky130_fd_sc_hd__conb_1 conb_T35Y52 (.HI(tie_high_T35Y52), .LO(tie_low_T35Y52));
  sky130_fd_sc_hd__conb_1 conb_T35Y53 (.HI(tie_high_T35Y53), .LO(tie_low_T35Y53));
  sky130_fd_sc_hd__conb_1 conb_T35Y54 (.HI(tie_high_T35Y54), .LO(tie_low_T35Y54));
  sky130_fd_sc_hd__conb_1 conb_T35Y55 (.HI(tie_high_T35Y55), .LO(tie_low_T35Y55));
  sky130_fd_sc_hd__conb_1 conb_T35Y56 (.HI(tie_high_T35Y56), .LO(tie_low_T35Y56));
  sky130_fd_sc_hd__conb_1 conb_T35Y57 (.HI(tie_high_T35Y57), .LO(tie_low_T35Y57));
  sky130_fd_sc_hd__conb_1 conb_T35Y58 (.HI(tie_high_T35Y58), .LO(tie_low_T35Y58));
  sky130_fd_sc_hd__conb_1 conb_T35Y59 (.HI(tie_high_T35Y59), .LO(tie_low_T35Y59));
  sky130_fd_sc_hd__conb_1 conb_T35Y6 (.HI(tie_high_T35Y6), .LO(tie_low_T35Y6));
  sky130_fd_sc_hd__conb_1 conb_T35Y60 (.HI(tie_high_T35Y60), .LO(tie_low_T35Y60));
  sky130_fd_sc_hd__conb_1 conb_T35Y61 (.HI(tie_high_T35Y61), .LO(tie_low_T35Y61));
  sky130_fd_sc_hd__conb_1 conb_T35Y62 (.HI(tie_high_T35Y62), .LO(tie_low_T35Y62));
  sky130_fd_sc_hd__conb_1 conb_T35Y63 (.HI(tie_high_T35Y63), .LO(tie_low_T35Y63));
  sky130_fd_sc_hd__conb_1 conb_T35Y64 (.HI(tie_high_T35Y64), .LO(tie_low_T35Y64));
  sky130_fd_sc_hd__conb_1 conb_T35Y65 (.HI(tie_high_T35Y65), .LO(tie_low_T35Y65));
  sky130_fd_sc_hd__conb_1 conb_T35Y66 (.HI(tie_high_T35Y66), .LO(tie_low_T35Y66));
  sky130_fd_sc_hd__conb_1 conb_T35Y67 (.HI(tie_high_T35Y67), .LO(tie_low_T35Y67));
  sky130_fd_sc_hd__conb_1 conb_T35Y68 (.HI(tie_high_T35Y68), .LO(tie_low_T35Y68));
  sky130_fd_sc_hd__conb_1 conb_T35Y69 (.HI(tie_high_T35Y69), .LO(tie_low_T35Y69));
  sky130_fd_sc_hd__conb_1 conb_T35Y7 (.HI(tie_high_T35Y7), .LO(tie_low_T35Y7));
  sky130_fd_sc_hd__conb_1 conb_T35Y70 (.HI(tie_high_T35Y70), .LO(tie_low_T35Y70));
  sky130_fd_sc_hd__conb_1 conb_T35Y71 (.HI(tie_high_T35Y71), .LO(tie_low_T35Y71));
  sky130_fd_sc_hd__conb_1 conb_T35Y72 (.HI(tie_high_T35Y72), .LO(tie_low_T35Y72));
  sky130_fd_sc_hd__conb_1 conb_T35Y73 (.HI(tie_high_T35Y73), .LO(tie_low_T35Y73));
  sky130_fd_sc_hd__conb_1 conb_T35Y74 (.HI(tie_high_T35Y74), .LO(tie_low_T35Y74));
  sky130_fd_sc_hd__conb_1 conb_T35Y75 (.HI(tie_high_T35Y75), .LO(tie_low_T35Y75));
  sky130_fd_sc_hd__conb_1 conb_T35Y76 (.HI(tie_high_T35Y76), .LO(tie_low_T35Y76));
  sky130_fd_sc_hd__conb_1 conb_T35Y77 (.HI(tie_high_T35Y77), .LO(tie_low_T35Y77));
  sky130_fd_sc_hd__conb_1 conb_T35Y78 (.HI(tie_high_T35Y78), .LO(tie_low_T35Y78));
  sky130_fd_sc_hd__conb_1 conb_T35Y79 (.HI(tie_high_T35Y79), .LO(tie_low_T35Y79));
  sky130_fd_sc_hd__conb_1 conb_T35Y8 (.HI(tie_high_T35Y8), .LO(tie_low_T35Y8));
  sky130_fd_sc_hd__conb_1 conb_T35Y80 (.HI(tie_high_T35Y80), .LO(tie_low_T35Y80));
  sky130_fd_sc_hd__conb_1 conb_T35Y81 (.HI(tie_high_T35Y81), .LO(tie_low_T35Y81));
  sky130_fd_sc_hd__conb_1 conb_T35Y82 (.HI(tie_high_T35Y82), .LO(tie_low_T35Y82));
  sky130_fd_sc_hd__conb_1 conb_T35Y83 (.HI(tie_high_T35Y83), .LO(tie_low_T35Y83));
  sky130_fd_sc_hd__conb_1 conb_T35Y84 (.HI(tie_high_T35Y84), .LO(tie_low_T35Y84));
  sky130_fd_sc_hd__conb_1 conb_T35Y85 (.HI(tie_high_T35Y85), .LO(tie_low_T35Y85));
  sky130_fd_sc_hd__conb_1 conb_T35Y86 (.HI(tie_high_T35Y86), .LO(tie_low_T35Y86));
  sky130_fd_sc_hd__conb_1 conb_T35Y87 (.HI(tie_high_T35Y87), .LO(tie_low_T35Y87));
  sky130_fd_sc_hd__conb_1 conb_T35Y88 (.HI(tie_high_T35Y88), .LO(tie_low_T35Y88));
  sky130_fd_sc_hd__conb_1 conb_T35Y89 (.HI(tie_high_T35Y89), .LO(tie_low_T35Y89));
  sky130_fd_sc_hd__conb_1 conb_T35Y9 (.HI(tie_high_T35Y9), .LO(tie_low_T35Y9));
  sky130_fd_sc_hd__conb_1 conb_T3Y0 (.HI(tie_high_T3Y0), .LO(tie_low_T3Y0));
  sky130_fd_sc_hd__conb_1 conb_T3Y1 (.HI(tie_high_T3Y1), .LO(tie_low_T3Y1));
  sky130_fd_sc_hd__conb_1 conb_T3Y10 (.HI(tie_high_T3Y10), .LO(tie_low_T3Y10));
  sky130_fd_sc_hd__conb_1 conb_T3Y11 (.HI(tie_high_T3Y11), .LO(tie_low_T3Y11));
  sky130_fd_sc_hd__conb_1 conb_T3Y12 (.HI(tie_high_T3Y12), .LO(tie_low_T3Y12));
  sky130_fd_sc_hd__conb_1 conb_T3Y13 (.HI(tie_high_T3Y13), .LO(tie_low_T3Y13));
  sky130_fd_sc_hd__conb_1 conb_T3Y14 (.HI(tie_high_T3Y14), .LO(tie_low_T3Y14));
  sky130_fd_sc_hd__conb_1 conb_T3Y15 (.HI(tie_high_T3Y15), .LO(tie_low_T3Y15));
  sky130_fd_sc_hd__conb_1 conb_T3Y16 (.HI(tie_high_T3Y16), .LO(tie_low_T3Y16));
  sky130_fd_sc_hd__conb_1 conb_T3Y17 (.HI(tie_high_T3Y17), .LO(tie_low_T3Y17));
  sky130_fd_sc_hd__conb_1 conb_T3Y18 (.HI(tie_high_T3Y18), .LO(tie_low_T3Y18));
  sky130_fd_sc_hd__conb_1 conb_T3Y19 (.HI(tie_high_T3Y19), .LO(tie_low_T3Y19));
  sky130_fd_sc_hd__conb_1 conb_T3Y2 (.HI(tie_high_T3Y2), .LO(tie_low_T3Y2));
  sky130_fd_sc_hd__conb_1 conb_T3Y20 (.HI(tie_high_T3Y20), .LO(tie_low_T3Y20));
  sky130_fd_sc_hd__conb_1 conb_T3Y21 (.HI(tie_high_T3Y21), .LO(tie_low_T3Y21));
  sky130_fd_sc_hd__conb_1 conb_T3Y22 (.HI(tie_high_T3Y22), .LO(tie_low_T3Y22));
  sky130_fd_sc_hd__conb_1 conb_T3Y23 (.HI(tie_high_T3Y23), .LO(tie_low_T3Y23));
  sky130_fd_sc_hd__conb_1 conb_T3Y24 (.HI(tie_high_T3Y24), .LO(tie_low_T3Y24));
  sky130_fd_sc_hd__conb_1 conb_T3Y25 (.HI(tie_high_T3Y25), .LO(tie_low_T3Y25));
  sky130_fd_sc_hd__conb_1 conb_T3Y26 (.HI(tie_high_T3Y26), .LO(tie_low_T3Y26));
  sky130_fd_sc_hd__conb_1 conb_T3Y27 (.HI(tie_high_T3Y27), .LO(tie_low_T3Y27));
  sky130_fd_sc_hd__conb_1 conb_T3Y28 (.HI(tie_high_T3Y28), .LO(tie_low_T3Y28));
  sky130_fd_sc_hd__conb_1 conb_T3Y29 (.HI(tie_high_T3Y29), .LO(tie_low_T3Y29));
  sky130_fd_sc_hd__conb_1 conb_T3Y3 (.HI(tie_high_T3Y3), .LO(tie_low_T3Y3));
  sky130_fd_sc_hd__conb_1 conb_T3Y30 (.HI(tie_high_T3Y30), .LO(tie_low_T3Y30));
  sky130_fd_sc_hd__conb_1 conb_T3Y31 (.HI(tie_high_T3Y31), .LO(tie_low_T3Y31));
  sky130_fd_sc_hd__conb_1 conb_T3Y32 (.HI(tie_high_T3Y32), .LO(tie_low_T3Y32));
  sky130_fd_sc_hd__conb_1 conb_T3Y33 (.HI(tie_high_T3Y33), .LO(tie_low_T3Y33));
  sky130_fd_sc_hd__conb_1 conb_T3Y34 (.HI(tie_high_T3Y34), .LO(tie_low_T3Y34));
  sky130_fd_sc_hd__conb_1 conb_T3Y35 (.HI(tie_high_T3Y35), .LO(tie_low_T3Y35));
  sky130_fd_sc_hd__conb_1 conb_T3Y36 (.HI(tie_high_T3Y36), .LO(tie_low_T3Y36));
  sky130_fd_sc_hd__conb_1 conb_T3Y37 (.HI(tie_high_T3Y37), .LO(tie_low_T3Y37));
  sky130_fd_sc_hd__conb_1 conb_T3Y38 (.HI(tie_high_T3Y38), .LO(tie_low_T3Y38));
  sky130_fd_sc_hd__conb_1 conb_T3Y39 (.HI(tie_high_T3Y39), .LO(tie_low_T3Y39));
  sky130_fd_sc_hd__conb_1 conb_T3Y4 (.HI(tie_high_T3Y4), .LO(tie_low_T3Y4));
  sky130_fd_sc_hd__conb_1 conb_T3Y40 (.HI(tie_high_T3Y40), .LO(tie_low_T3Y40));
  sky130_fd_sc_hd__conb_1 conb_T3Y41 (.HI(tie_high_T3Y41), .LO(tie_low_T3Y41));
  sky130_fd_sc_hd__conb_1 conb_T3Y42 (.HI(tie_high_T3Y42), .LO(tie_low_T3Y42));
  sky130_fd_sc_hd__conb_1 conb_T3Y43 (.HI(tie_high_T3Y43), .LO(tie_low_T3Y43));
  sky130_fd_sc_hd__conb_1 conb_T3Y44 (.HI(tie_high_T3Y44), .LO(tie_low_T3Y44));
  sky130_fd_sc_hd__conb_1 conb_T3Y45 (.HI(tie_high_T3Y45), .LO(tie_low_T3Y45));
  sky130_fd_sc_hd__conb_1 conb_T3Y46 (.HI(tie_high_T3Y46), .LO(tie_low_T3Y46));
  sky130_fd_sc_hd__conb_1 conb_T3Y47 (.HI(tie_high_T3Y47), .LO(tie_low_T3Y47));
  sky130_fd_sc_hd__conb_1 conb_T3Y48 (.HI(tie_high_T3Y48), .LO(tie_low_T3Y48));
  sky130_fd_sc_hd__conb_1 conb_T3Y49 (.HI(tie_high_T3Y49), .LO(tie_low_T3Y49));
  sky130_fd_sc_hd__conb_1 conb_T3Y5 (.HI(tie_high_T3Y5), .LO(tie_low_T3Y5));
  sky130_fd_sc_hd__conb_1 conb_T3Y50 (.HI(tie_high_T3Y50), .LO(tie_low_T3Y50));
  sky130_fd_sc_hd__conb_1 conb_T3Y51 (.HI(tie_high_T3Y51), .LO(tie_low_T3Y51));
  sky130_fd_sc_hd__conb_1 conb_T3Y52 (.HI(tie_high_T3Y52), .LO(tie_low_T3Y52));
  sky130_fd_sc_hd__conb_1 conb_T3Y53 (.HI(tie_high_T3Y53), .LO(tie_low_T3Y53));
  sky130_fd_sc_hd__conb_1 conb_T3Y54 (.HI(tie_high_T3Y54), .LO(tie_low_T3Y54));
  sky130_fd_sc_hd__conb_1 conb_T3Y55 (.HI(tie_high_T3Y55), .LO(tie_low_T3Y55));
  sky130_fd_sc_hd__conb_1 conb_T3Y56 (.HI(tie_high_T3Y56), .LO(tie_low_T3Y56));
  sky130_fd_sc_hd__conb_1 conb_T3Y57 (.HI(tie_high_T3Y57), .LO(tie_low_T3Y57));
  sky130_fd_sc_hd__conb_1 conb_T3Y58 (.HI(tie_high_T3Y58), .LO(tie_low_T3Y58));
  sky130_fd_sc_hd__conb_1 conb_T3Y59 (.HI(tie_high_T3Y59), .LO(tie_low_T3Y59));
  sky130_fd_sc_hd__conb_1 conb_T3Y6 (.HI(tie_high_T3Y6), .LO(tie_low_T3Y6));
  sky130_fd_sc_hd__conb_1 conb_T3Y60 (.HI(tie_high_T3Y60), .LO(tie_low_T3Y60));
  sky130_fd_sc_hd__conb_1 conb_T3Y61 (.HI(tie_high_T3Y61), .LO(tie_low_T3Y61));
  sky130_fd_sc_hd__conb_1 conb_T3Y62 (.HI(tie_high_T3Y62), .LO(tie_low_T3Y62));
  sky130_fd_sc_hd__conb_1 conb_T3Y63 (.HI(tie_high_T3Y63), .LO(tie_low_T3Y63));
  sky130_fd_sc_hd__conb_1 conb_T3Y64 (.HI(tie_high_T3Y64), .LO(tie_low_T3Y64));
  sky130_fd_sc_hd__conb_1 conb_T3Y65 (.HI(tie_high_T3Y65), .LO(tie_low_T3Y65));
  sky130_fd_sc_hd__conb_1 conb_T3Y66 (.HI(tie_high_T3Y66), .LO(tie_low_T3Y66));
  sky130_fd_sc_hd__conb_1 conb_T3Y67 (.HI(tie_high_T3Y67), .LO(tie_low_T3Y67));
  sky130_fd_sc_hd__conb_1 conb_T3Y68 (.HI(tie_high_T3Y68), .LO(tie_low_T3Y68));
  sky130_fd_sc_hd__conb_1 conb_T3Y69 (.HI(tie_high_T3Y69), .LO(tie_low_T3Y69));
  sky130_fd_sc_hd__conb_1 conb_T3Y7 (.HI(tie_high_T3Y7), .LO(tie_low_T3Y7));
  sky130_fd_sc_hd__conb_1 conb_T3Y70 (.HI(tie_high_T3Y70), .LO(tie_low_T3Y70));
  sky130_fd_sc_hd__conb_1 conb_T3Y71 (.HI(tie_high_T3Y71), .LO(tie_low_T3Y71));
  sky130_fd_sc_hd__conb_1 conb_T3Y72 (.HI(tie_high_T3Y72), .LO(tie_low_T3Y72));
  sky130_fd_sc_hd__conb_1 conb_T3Y73 (.HI(tie_high_T3Y73), .LO(tie_low_T3Y73));
  sky130_fd_sc_hd__conb_1 conb_T3Y74 (.HI(tie_high_T3Y74), .LO(tie_low_T3Y74));
  sky130_fd_sc_hd__conb_1 conb_T3Y75 (.HI(tie_high_T3Y75), .LO(tie_low_T3Y75));
  sky130_fd_sc_hd__conb_1 conb_T3Y76 (.HI(tie_high_T3Y76), .LO(tie_low_T3Y76));
  sky130_fd_sc_hd__conb_1 conb_T3Y77 (.HI(tie_high_T3Y77), .LO(tie_low_T3Y77));
  sky130_fd_sc_hd__conb_1 conb_T3Y78 (.HI(tie_high_T3Y78), .LO(tie_low_T3Y78));
  sky130_fd_sc_hd__conb_1 conb_T3Y79 (.HI(tie_high_T3Y79), .LO(tie_low_T3Y79));
  sky130_fd_sc_hd__conb_1 conb_T3Y8 (.HI(tie_high_T3Y8), .LO(tie_low_T3Y8));
  sky130_fd_sc_hd__conb_1 conb_T3Y80 (.HI(tie_high_T3Y80), .LO(tie_low_T3Y80));
  sky130_fd_sc_hd__conb_1 conb_T3Y81 (.HI(tie_high_T3Y81), .LO(tie_low_T3Y81));
  sky130_fd_sc_hd__conb_1 conb_T3Y82 (.HI(tie_high_T3Y82), .LO(tie_low_T3Y82));
  sky130_fd_sc_hd__conb_1 conb_T3Y83 (.HI(tie_high_T3Y83), .LO(tie_low_T3Y83));
  sky130_fd_sc_hd__conb_1 conb_T3Y84 (.HI(tie_high_T3Y84), .LO(tie_low_T3Y84));
  sky130_fd_sc_hd__conb_1 conb_T3Y85 (.HI(tie_high_T3Y85), .LO(tie_low_T3Y85));
  sky130_fd_sc_hd__conb_1 conb_T3Y86 (.HI(tie_high_T3Y86), .LO(tie_low_T3Y86));
  sky130_fd_sc_hd__conb_1 conb_T3Y87 (.HI(tie_high_T3Y87), .LO(tie_low_T3Y87));
  sky130_fd_sc_hd__conb_1 conb_T3Y88 (.HI(tie_high_T3Y88), .LO(tie_low_T3Y88));
  sky130_fd_sc_hd__conb_1 conb_T3Y89 (.HI(tie_high_T3Y89), .LO(tie_low_T3Y89));
  sky130_fd_sc_hd__conb_1 conb_T3Y9 (.HI(tie_high_T3Y9), .LO(tie_low_T3Y9));
  sky130_fd_sc_hd__conb_1 conb_T4Y0 (.HI(tie_high_T4Y0), .LO(tie_low_T4Y0));
  sky130_fd_sc_hd__conb_1 conb_T4Y1 (.HI(tie_high_T4Y1), .LO(tie_low_T4Y1));
  sky130_fd_sc_hd__conb_1 conb_T4Y10 (.HI(tie_high_T4Y10), .LO(tie_low_T4Y10));
  sky130_fd_sc_hd__conb_1 conb_T4Y11 (.HI(tie_high_T4Y11), .LO(tie_low_T4Y11));
  sky130_fd_sc_hd__conb_1 conb_T4Y12 (.HI(tie_high_T4Y12), .LO(tie_low_T4Y12));
  sky130_fd_sc_hd__conb_1 conb_T4Y13 (.HI(tie_high_T4Y13), .LO(tie_low_T4Y13));
  sky130_fd_sc_hd__conb_1 conb_T4Y14 (.HI(tie_high_T4Y14), .LO(tie_low_T4Y14));
  sky130_fd_sc_hd__conb_1 conb_T4Y15 (.HI(tie_high_T4Y15), .LO(tie_low_T4Y15));
  sky130_fd_sc_hd__conb_1 conb_T4Y16 (.HI(tie_high_T4Y16), .LO(tie_low_T4Y16));
  sky130_fd_sc_hd__conb_1 conb_T4Y17 (.HI(tie_high_T4Y17), .LO(tie_low_T4Y17));
  sky130_fd_sc_hd__conb_1 conb_T4Y18 (.HI(tie_high_T4Y18), .LO(tie_low_T4Y18));
  sky130_fd_sc_hd__conb_1 conb_T4Y19 (.HI(tie_high_T4Y19), .LO(tie_low_T4Y19));
  sky130_fd_sc_hd__conb_1 conb_T4Y2 (.HI(tie_high_T4Y2), .LO(tie_low_T4Y2));
  sky130_fd_sc_hd__conb_1 conb_T4Y20 (.HI(tie_high_T4Y20), .LO(tie_low_T4Y20));
  sky130_fd_sc_hd__conb_1 conb_T4Y21 (.HI(tie_high_T4Y21), .LO(tie_low_T4Y21));
  sky130_fd_sc_hd__conb_1 conb_T4Y22 (.HI(tie_high_T4Y22), .LO(tie_low_T4Y22));
  sky130_fd_sc_hd__conb_1 conb_T4Y23 (.HI(tie_high_T4Y23), .LO(tie_low_T4Y23));
  sky130_fd_sc_hd__conb_1 conb_T4Y24 (.HI(tie_high_T4Y24), .LO(tie_low_T4Y24));
  sky130_fd_sc_hd__conb_1 conb_T4Y25 (.HI(tie_high_T4Y25), .LO(tie_low_T4Y25));
  sky130_fd_sc_hd__conb_1 conb_T4Y26 (.HI(tie_high_T4Y26), .LO(tie_low_T4Y26));
  sky130_fd_sc_hd__conb_1 conb_T4Y27 (.HI(tie_high_T4Y27), .LO(tie_low_T4Y27));
  sky130_fd_sc_hd__conb_1 conb_T4Y28 (.HI(tie_high_T4Y28), .LO(tie_low_T4Y28));
  sky130_fd_sc_hd__conb_1 conb_T4Y29 (.HI(tie_high_T4Y29), .LO(tie_low_T4Y29));
  sky130_fd_sc_hd__conb_1 conb_T4Y3 (.HI(tie_high_T4Y3), .LO(tie_low_T4Y3));
  sky130_fd_sc_hd__conb_1 conb_T4Y30 (.HI(tie_high_T4Y30), .LO(tie_low_T4Y30));
  sky130_fd_sc_hd__conb_1 conb_T4Y31 (.HI(tie_high_T4Y31), .LO(tie_low_T4Y31));
  sky130_fd_sc_hd__conb_1 conb_T4Y32 (.HI(tie_high_T4Y32), .LO(tie_low_T4Y32));
  sky130_fd_sc_hd__conb_1 conb_T4Y33 (.HI(tie_high_T4Y33), .LO(tie_low_T4Y33));
  sky130_fd_sc_hd__conb_1 conb_T4Y34 (.HI(tie_high_T4Y34), .LO(tie_low_T4Y34));
  sky130_fd_sc_hd__conb_1 conb_T4Y35 (.HI(tie_high_T4Y35), .LO(tie_low_T4Y35));
  sky130_fd_sc_hd__conb_1 conb_T4Y36 (.HI(tie_high_T4Y36), .LO(tie_low_T4Y36));
  sky130_fd_sc_hd__conb_1 conb_T4Y37 (.HI(tie_high_T4Y37), .LO(tie_low_T4Y37));
  sky130_fd_sc_hd__conb_1 conb_T4Y38 (.HI(tie_high_T4Y38), .LO(tie_low_T4Y38));
  sky130_fd_sc_hd__conb_1 conb_T4Y39 (.HI(tie_high_T4Y39), .LO(tie_low_T4Y39));
  sky130_fd_sc_hd__conb_1 conb_T4Y4 (.HI(tie_high_T4Y4), .LO(tie_low_T4Y4));
  sky130_fd_sc_hd__conb_1 conb_T4Y40 (.HI(tie_high_T4Y40), .LO(tie_low_T4Y40));
  sky130_fd_sc_hd__conb_1 conb_T4Y41 (.HI(tie_high_T4Y41), .LO(tie_low_T4Y41));
  sky130_fd_sc_hd__conb_1 conb_T4Y42 (.HI(tie_high_T4Y42), .LO(tie_low_T4Y42));
  sky130_fd_sc_hd__conb_1 conb_T4Y43 (.HI(tie_high_T4Y43), .LO(tie_low_T4Y43));
  sky130_fd_sc_hd__conb_1 conb_T4Y44 (.HI(tie_high_T4Y44), .LO(tie_low_T4Y44));
  sky130_fd_sc_hd__conb_1 conb_T4Y45 (.HI(tie_high_T4Y45), .LO(tie_low_T4Y45));
  sky130_fd_sc_hd__conb_1 conb_T4Y46 (.HI(tie_high_T4Y46), .LO(tie_low_T4Y46));
  sky130_fd_sc_hd__conb_1 conb_T4Y47 (.HI(tie_high_T4Y47), .LO(tie_low_T4Y47));
  sky130_fd_sc_hd__conb_1 conb_T4Y48 (.HI(tie_high_T4Y48), .LO(tie_low_T4Y48));
  sky130_fd_sc_hd__conb_1 conb_T4Y49 (.HI(tie_high_T4Y49), .LO(tie_low_T4Y49));
  sky130_fd_sc_hd__conb_1 conb_T4Y5 (.HI(tie_high_T4Y5), .LO(tie_low_T4Y5));
  sky130_fd_sc_hd__conb_1 conb_T4Y50 (.HI(tie_high_T4Y50), .LO(tie_low_T4Y50));
  sky130_fd_sc_hd__conb_1 conb_T4Y51 (.HI(tie_high_T4Y51), .LO(tie_low_T4Y51));
  sky130_fd_sc_hd__conb_1 conb_T4Y52 (.HI(tie_high_T4Y52), .LO(tie_low_T4Y52));
  sky130_fd_sc_hd__conb_1 conb_T4Y53 (.HI(tie_high_T4Y53), .LO(tie_low_T4Y53));
  sky130_fd_sc_hd__conb_1 conb_T4Y54 (.HI(tie_high_T4Y54), .LO(tie_low_T4Y54));
  sky130_fd_sc_hd__conb_1 conb_T4Y55 (.HI(tie_high_T4Y55), .LO(tie_low_T4Y55));
  sky130_fd_sc_hd__conb_1 conb_T4Y56 (.HI(tie_high_T4Y56), .LO(tie_low_T4Y56));
  sky130_fd_sc_hd__conb_1 conb_T4Y57 (.HI(tie_high_T4Y57), .LO(tie_low_T4Y57));
  sky130_fd_sc_hd__conb_1 conb_T4Y58 (.HI(tie_high_T4Y58), .LO(tie_low_T4Y58));
  sky130_fd_sc_hd__conb_1 conb_T4Y59 (.HI(tie_high_T4Y59), .LO(tie_low_T4Y59));
  sky130_fd_sc_hd__conb_1 conb_T4Y6 (.HI(tie_high_T4Y6), .LO(tie_low_T4Y6));
  sky130_fd_sc_hd__conb_1 conb_T4Y60 (.HI(tie_high_T4Y60), .LO(tie_low_T4Y60));
  sky130_fd_sc_hd__conb_1 conb_T4Y61 (.HI(tie_high_T4Y61), .LO(tie_low_T4Y61));
  sky130_fd_sc_hd__conb_1 conb_T4Y62 (.HI(tie_high_T4Y62), .LO(tie_low_T4Y62));
  sky130_fd_sc_hd__conb_1 conb_T4Y63 (.HI(tie_high_T4Y63), .LO(tie_low_T4Y63));
  sky130_fd_sc_hd__conb_1 conb_T4Y64 (.HI(tie_high_T4Y64), .LO(tie_low_T4Y64));
  sky130_fd_sc_hd__conb_1 conb_T4Y65 (.HI(tie_high_T4Y65), .LO(tie_low_T4Y65));
  sky130_fd_sc_hd__conb_1 conb_T4Y66 (.HI(tie_high_T4Y66), .LO(tie_low_T4Y66));
  sky130_fd_sc_hd__conb_1 conb_T4Y67 (.HI(tie_high_T4Y67), .LO(tie_low_T4Y67));
  sky130_fd_sc_hd__conb_1 conb_T4Y68 (.HI(tie_high_T4Y68), .LO(tie_low_T4Y68));
  sky130_fd_sc_hd__conb_1 conb_T4Y69 (.HI(tie_high_T4Y69), .LO(tie_low_T4Y69));
  sky130_fd_sc_hd__conb_1 conb_T4Y7 (.HI(tie_high_T4Y7), .LO(tie_low_T4Y7));
  sky130_fd_sc_hd__conb_1 conb_T4Y70 (.HI(tie_high_T4Y70), .LO(tie_low_T4Y70));
  sky130_fd_sc_hd__conb_1 conb_T4Y71 (.HI(tie_high_T4Y71), .LO(tie_low_T4Y71));
  sky130_fd_sc_hd__conb_1 conb_T4Y72 (.HI(tie_high_T4Y72), .LO(tie_low_T4Y72));
  sky130_fd_sc_hd__conb_1 conb_T4Y73 (.HI(tie_high_T4Y73), .LO(tie_low_T4Y73));
  sky130_fd_sc_hd__conb_1 conb_T4Y74 (.HI(tie_high_T4Y74), .LO(tie_low_T4Y74));
  sky130_fd_sc_hd__conb_1 conb_T4Y75 (.HI(tie_high_T4Y75), .LO(tie_low_T4Y75));
  sky130_fd_sc_hd__conb_1 conb_T4Y76 (.HI(tie_high_T4Y76), .LO(tie_low_T4Y76));
  sky130_fd_sc_hd__conb_1 conb_T4Y77 (.HI(tie_high_T4Y77), .LO(tie_low_T4Y77));
  sky130_fd_sc_hd__conb_1 conb_T4Y78 (.HI(tie_high_T4Y78), .LO(tie_low_T4Y78));
  sky130_fd_sc_hd__conb_1 conb_T4Y79 (.HI(tie_high_T4Y79), .LO(tie_low_T4Y79));
  sky130_fd_sc_hd__conb_1 conb_T4Y8 (.HI(tie_high_T4Y8), .LO(tie_low_T4Y8));
  sky130_fd_sc_hd__conb_1 conb_T4Y80 (.HI(tie_high_T4Y80), .LO(tie_low_T4Y80));
  sky130_fd_sc_hd__conb_1 conb_T4Y81 (.HI(tie_high_T4Y81), .LO(tie_low_T4Y81));
  sky130_fd_sc_hd__conb_1 conb_T4Y82 (.HI(tie_high_T4Y82), .LO(tie_low_T4Y82));
  sky130_fd_sc_hd__conb_1 conb_T4Y83 (.HI(tie_high_T4Y83), .LO(tie_low_T4Y83));
  sky130_fd_sc_hd__conb_1 conb_T4Y84 (.HI(tie_high_T4Y84), .LO(tie_low_T4Y84));
  sky130_fd_sc_hd__conb_1 conb_T4Y85 (.HI(tie_high_T4Y85), .LO(tie_low_T4Y85));
  sky130_fd_sc_hd__conb_1 conb_T4Y86 (.HI(tie_high_T4Y86), .LO(tie_low_T4Y86));
  sky130_fd_sc_hd__conb_1 conb_T4Y87 (.HI(tie_high_T4Y87), .LO(tie_low_T4Y87));
  sky130_fd_sc_hd__conb_1 conb_T4Y88 (.HI(tie_high_T4Y88), .LO(tie_low_T4Y88));
  sky130_fd_sc_hd__conb_1 conb_T4Y89 (.HI(tie_high_T4Y89), .LO(tie_low_T4Y89));
  sky130_fd_sc_hd__conb_1 conb_T4Y9 (.HI(tie_high_T4Y9), .LO(tie_low_T4Y9));
  sky130_fd_sc_hd__conb_1 conb_T5Y0 (.HI(tie_high_T5Y0), .LO(tie_low_T5Y0));
  sky130_fd_sc_hd__conb_1 conb_T5Y1 (.HI(tie_high_T5Y1), .LO(tie_low_T5Y1));
  sky130_fd_sc_hd__conb_1 conb_T5Y10 (.HI(tie_high_T5Y10), .LO(tie_low_T5Y10));
  sky130_fd_sc_hd__conb_1 conb_T5Y11 (.HI(tie_high_T5Y11), .LO(tie_low_T5Y11));
  sky130_fd_sc_hd__conb_1 conb_T5Y12 (.HI(tie_high_T5Y12), .LO(tie_low_T5Y12));
  sky130_fd_sc_hd__conb_1 conb_T5Y13 (.HI(tie_high_T5Y13), .LO(tie_low_T5Y13));
  sky130_fd_sc_hd__conb_1 conb_T5Y14 (.HI(tie_high_T5Y14), .LO(tie_low_T5Y14));
  sky130_fd_sc_hd__conb_1 conb_T5Y15 (.HI(tie_high_T5Y15), .LO(tie_low_T5Y15));
  sky130_fd_sc_hd__conb_1 conb_T5Y16 (.HI(tie_high_T5Y16), .LO(tie_low_T5Y16));
  sky130_fd_sc_hd__conb_1 conb_T5Y17 (.HI(tie_high_T5Y17), .LO(tie_low_T5Y17));
  sky130_fd_sc_hd__conb_1 conb_T5Y18 (.HI(tie_high_T5Y18), .LO(tie_low_T5Y18));
  sky130_fd_sc_hd__conb_1 conb_T5Y19 (.HI(tie_high_T5Y19), .LO(tie_low_T5Y19));
  sky130_fd_sc_hd__conb_1 conb_T5Y2 (.HI(tie_high_T5Y2), .LO(tie_low_T5Y2));
  sky130_fd_sc_hd__conb_1 conb_T5Y20 (.HI(tie_high_T5Y20), .LO(tie_low_T5Y20));
  sky130_fd_sc_hd__conb_1 conb_T5Y21 (.HI(tie_high_T5Y21), .LO(tie_low_T5Y21));
  sky130_fd_sc_hd__conb_1 conb_T5Y22 (.HI(tie_high_T5Y22), .LO(tie_low_T5Y22));
  sky130_fd_sc_hd__conb_1 conb_T5Y23 (.HI(tie_high_T5Y23), .LO(tie_low_T5Y23));
  sky130_fd_sc_hd__conb_1 conb_T5Y24 (.HI(tie_high_T5Y24), .LO(tie_low_T5Y24));
  sky130_fd_sc_hd__conb_1 conb_T5Y25 (.HI(tie_high_T5Y25), .LO(tie_low_T5Y25));
  sky130_fd_sc_hd__conb_1 conb_T5Y26 (.HI(tie_high_T5Y26), .LO(tie_low_T5Y26));
  sky130_fd_sc_hd__conb_1 conb_T5Y27 (.HI(tie_high_T5Y27), .LO(tie_low_T5Y27));
  sky130_fd_sc_hd__conb_1 conb_T5Y28 (.HI(tie_high_T5Y28), .LO(tie_low_T5Y28));
  sky130_fd_sc_hd__conb_1 conb_T5Y29 (.HI(tie_high_T5Y29), .LO(tie_low_T5Y29));
  sky130_fd_sc_hd__conb_1 conb_T5Y3 (.HI(tie_high_T5Y3), .LO(tie_low_T5Y3));
  sky130_fd_sc_hd__conb_1 conb_T5Y30 (.HI(tie_high_T5Y30), .LO(tie_low_T5Y30));
  sky130_fd_sc_hd__conb_1 conb_T5Y31 (.HI(tie_high_T5Y31), .LO(tie_low_T5Y31));
  sky130_fd_sc_hd__conb_1 conb_T5Y32 (.HI(tie_high_T5Y32), .LO(tie_low_T5Y32));
  sky130_fd_sc_hd__conb_1 conb_T5Y33 (.HI(tie_high_T5Y33), .LO(tie_low_T5Y33));
  sky130_fd_sc_hd__conb_1 conb_T5Y34 (.HI(tie_high_T5Y34), .LO(tie_low_T5Y34));
  sky130_fd_sc_hd__conb_1 conb_T5Y35 (.HI(tie_high_T5Y35), .LO(tie_low_T5Y35));
  sky130_fd_sc_hd__conb_1 conb_T5Y36 (.HI(tie_high_T5Y36), .LO(tie_low_T5Y36));
  sky130_fd_sc_hd__conb_1 conb_T5Y37 (.HI(tie_high_T5Y37), .LO(tie_low_T5Y37));
  sky130_fd_sc_hd__conb_1 conb_T5Y38 (.HI(tie_high_T5Y38), .LO(tie_low_T5Y38));
  sky130_fd_sc_hd__conb_1 conb_T5Y39 (.HI(tie_high_T5Y39), .LO(tie_low_T5Y39));
  sky130_fd_sc_hd__conb_1 conb_T5Y4 (.HI(tie_high_T5Y4), .LO(tie_low_T5Y4));
  sky130_fd_sc_hd__conb_1 conb_T5Y40 (.HI(tie_high_T5Y40), .LO(tie_low_T5Y40));
  sky130_fd_sc_hd__conb_1 conb_T5Y41 (.HI(tie_high_T5Y41), .LO(tie_low_T5Y41));
  sky130_fd_sc_hd__conb_1 conb_T5Y42 (.HI(tie_high_T5Y42), .LO(tie_low_T5Y42));
  sky130_fd_sc_hd__conb_1 conb_T5Y43 (.HI(tie_high_T5Y43), .LO(tie_low_T5Y43));
  sky130_fd_sc_hd__conb_1 conb_T5Y44 (.HI(tie_high_T5Y44), .LO(tie_low_T5Y44));
  sky130_fd_sc_hd__conb_1 conb_T5Y45 (.HI(tie_high_T5Y45), .LO(tie_low_T5Y45));
  sky130_fd_sc_hd__conb_1 conb_T5Y46 (.HI(tie_high_T5Y46), .LO(tie_low_T5Y46));
  sky130_fd_sc_hd__conb_1 conb_T5Y47 (.HI(tie_high_T5Y47), .LO(tie_low_T5Y47));
  sky130_fd_sc_hd__conb_1 conb_T5Y48 (.HI(tie_high_T5Y48), .LO(tie_low_T5Y48));
  sky130_fd_sc_hd__conb_1 conb_T5Y49 (.HI(tie_high_T5Y49), .LO(tie_low_T5Y49));
  sky130_fd_sc_hd__conb_1 conb_T5Y5 (.HI(tie_high_T5Y5), .LO(tie_low_T5Y5));
  sky130_fd_sc_hd__conb_1 conb_T5Y50 (.HI(tie_high_T5Y50), .LO(tie_low_T5Y50));
  sky130_fd_sc_hd__conb_1 conb_T5Y51 (.HI(tie_high_T5Y51), .LO(tie_low_T5Y51));
  sky130_fd_sc_hd__conb_1 conb_T5Y52 (.HI(tie_high_T5Y52), .LO(tie_low_T5Y52));
  sky130_fd_sc_hd__conb_1 conb_T5Y53 (.HI(tie_high_T5Y53), .LO(tie_low_T5Y53));
  sky130_fd_sc_hd__conb_1 conb_T5Y54 (.HI(tie_high_T5Y54), .LO(tie_low_T5Y54));
  sky130_fd_sc_hd__conb_1 conb_T5Y55 (.HI(tie_high_T5Y55), .LO(tie_low_T5Y55));
  sky130_fd_sc_hd__conb_1 conb_T5Y56 (.HI(tie_high_T5Y56), .LO(tie_low_T5Y56));
  sky130_fd_sc_hd__conb_1 conb_T5Y57 (.HI(tie_high_T5Y57), .LO(tie_low_T5Y57));
  sky130_fd_sc_hd__conb_1 conb_T5Y58 (.HI(tie_high_T5Y58), .LO(tie_low_T5Y58));
  sky130_fd_sc_hd__conb_1 conb_T5Y59 (.HI(tie_high_T5Y59), .LO(tie_low_T5Y59));
  sky130_fd_sc_hd__conb_1 conb_T5Y6 (.HI(tie_high_T5Y6), .LO(tie_low_T5Y6));
  sky130_fd_sc_hd__conb_1 conb_T5Y60 (.HI(tie_high_T5Y60), .LO(tie_low_T5Y60));
  sky130_fd_sc_hd__conb_1 conb_T5Y61 (.HI(tie_high_T5Y61), .LO(tie_low_T5Y61));
  sky130_fd_sc_hd__conb_1 conb_T5Y62 (.HI(tie_high_T5Y62), .LO(tie_low_T5Y62));
  sky130_fd_sc_hd__conb_1 conb_T5Y63 (.HI(tie_high_T5Y63), .LO(tie_low_T5Y63));
  sky130_fd_sc_hd__conb_1 conb_T5Y64 (.HI(tie_high_T5Y64), .LO(tie_low_T5Y64));
  sky130_fd_sc_hd__conb_1 conb_T5Y65 (.HI(tie_high_T5Y65), .LO(tie_low_T5Y65));
  sky130_fd_sc_hd__conb_1 conb_T5Y66 (.HI(tie_high_T5Y66), .LO(tie_low_T5Y66));
  sky130_fd_sc_hd__conb_1 conb_T5Y67 (.HI(tie_high_T5Y67), .LO(tie_low_T5Y67));
  sky130_fd_sc_hd__conb_1 conb_T5Y68 (.HI(tie_high_T5Y68), .LO(tie_low_T5Y68));
  sky130_fd_sc_hd__conb_1 conb_T5Y69 (.HI(tie_high_T5Y69), .LO(tie_low_T5Y69));
  sky130_fd_sc_hd__conb_1 conb_T5Y7 (.HI(tie_high_T5Y7), .LO(tie_low_T5Y7));
  sky130_fd_sc_hd__conb_1 conb_T5Y70 (.HI(tie_high_T5Y70), .LO(tie_low_T5Y70));
  sky130_fd_sc_hd__conb_1 conb_T5Y71 (.HI(tie_high_T5Y71), .LO(tie_low_T5Y71));
  sky130_fd_sc_hd__conb_1 conb_T5Y72 (.HI(tie_high_T5Y72), .LO(tie_low_T5Y72));
  sky130_fd_sc_hd__conb_1 conb_T5Y73 (.HI(tie_high_T5Y73), .LO(tie_low_T5Y73));
  sky130_fd_sc_hd__conb_1 conb_T5Y74 (.HI(tie_high_T5Y74), .LO(tie_low_T5Y74));
  sky130_fd_sc_hd__conb_1 conb_T5Y75 (.HI(tie_high_T5Y75), .LO(tie_low_T5Y75));
  sky130_fd_sc_hd__conb_1 conb_T5Y76 (.HI(tie_high_T5Y76), .LO(tie_low_T5Y76));
  sky130_fd_sc_hd__conb_1 conb_T5Y77 (.HI(tie_high_T5Y77), .LO(tie_low_T5Y77));
  sky130_fd_sc_hd__conb_1 conb_T5Y78 (.HI(tie_high_T5Y78), .LO(tie_low_T5Y78));
  sky130_fd_sc_hd__conb_1 conb_T5Y79 (.HI(tie_high_T5Y79), .LO(tie_low_T5Y79));
  sky130_fd_sc_hd__conb_1 conb_T5Y8 (.HI(tie_high_T5Y8), .LO(tie_low_T5Y8));
  sky130_fd_sc_hd__conb_1 conb_T5Y80 (.HI(tie_high_T5Y80), .LO(tie_low_T5Y80));
  sky130_fd_sc_hd__conb_1 conb_T5Y81 (.HI(tie_high_T5Y81), .LO(tie_low_T5Y81));
  sky130_fd_sc_hd__conb_1 conb_T5Y82 (.HI(tie_high_T5Y82), .LO(tie_low_T5Y82));
  sky130_fd_sc_hd__conb_1 conb_T5Y83 (.HI(tie_high_T5Y83), .LO(tie_low_T5Y83));
  sky130_fd_sc_hd__conb_1 conb_T5Y84 (.HI(tie_high_T5Y84), .LO(tie_low_T5Y84));
  sky130_fd_sc_hd__conb_1 conb_T5Y85 (.HI(tie_high_T5Y85), .LO(tie_low_T5Y85));
  sky130_fd_sc_hd__conb_1 conb_T5Y86 (.HI(tie_high_T5Y86), .LO(tie_low_T5Y86));
  sky130_fd_sc_hd__conb_1 conb_T5Y87 (.HI(tie_high_T5Y87), .LO(tie_low_T5Y87));
  sky130_fd_sc_hd__conb_1 conb_T5Y88 (.HI(tie_high_T5Y88), .LO(tie_low_T5Y88));
  sky130_fd_sc_hd__conb_1 conb_T5Y89 (.HI(tie_high_T5Y89), .LO(tie_low_T5Y89));
  sky130_fd_sc_hd__conb_1 conb_T5Y9 (.HI(tie_high_T5Y9), .LO(tie_low_T5Y9));
  sky130_fd_sc_hd__conb_1 conb_T6Y0 (.HI(tie_high_T6Y0), .LO(tie_low_T6Y0));
  sky130_fd_sc_hd__conb_1 conb_T6Y1 (.HI(tie_high_T6Y1), .LO(tie_low_T6Y1));
  sky130_fd_sc_hd__conb_1 conb_T6Y10 (.HI(tie_high_T6Y10), .LO(tie_low_T6Y10));
  sky130_fd_sc_hd__conb_1 conb_T6Y11 (.HI(tie_high_T6Y11), .LO(tie_low_T6Y11));
  sky130_fd_sc_hd__conb_1 conb_T6Y12 (.HI(tie_high_T6Y12), .LO(tie_low_T6Y12));
  sky130_fd_sc_hd__conb_1 conb_T6Y13 (.HI(tie_high_T6Y13), .LO(tie_low_T6Y13));
  sky130_fd_sc_hd__conb_1 conb_T6Y14 (.HI(tie_high_T6Y14), .LO(tie_low_T6Y14));
  sky130_fd_sc_hd__conb_1 conb_T6Y15 (.HI(tie_high_T6Y15), .LO(tie_low_T6Y15));
  sky130_fd_sc_hd__conb_1 conb_T6Y16 (.HI(tie_high_T6Y16), .LO(tie_low_T6Y16));
  sky130_fd_sc_hd__conb_1 conb_T6Y17 (.HI(tie_high_T6Y17), .LO(tie_low_T6Y17));
  sky130_fd_sc_hd__conb_1 conb_T6Y18 (.HI(tie_high_T6Y18), .LO(tie_low_T6Y18));
  sky130_fd_sc_hd__conb_1 conb_T6Y19 (.HI(tie_high_T6Y19), .LO(tie_low_T6Y19));
  sky130_fd_sc_hd__conb_1 conb_T6Y2 (.HI(tie_high_T6Y2), .LO(tie_low_T6Y2));
  sky130_fd_sc_hd__conb_1 conb_T6Y20 (.HI(tie_high_T6Y20), .LO(tie_low_T6Y20));
  sky130_fd_sc_hd__conb_1 conb_T6Y21 (.HI(tie_high_T6Y21), .LO(tie_low_T6Y21));
  sky130_fd_sc_hd__conb_1 conb_T6Y22 (.HI(tie_high_T6Y22), .LO(tie_low_T6Y22));
  sky130_fd_sc_hd__conb_1 conb_T6Y23 (.HI(tie_high_T6Y23), .LO(tie_low_T6Y23));
  sky130_fd_sc_hd__conb_1 conb_T6Y24 (.HI(tie_high_T6Y24), .LO(tie_low_T6Y24));
  sky130_fd_sc_hd__conb_1 conb_T6Y25 (.HI(tie_high_T6Y25), .LO(tie_low_T6Y25));
  sky130_fd_sc_hd__conb_1 conb_T6Y26 (.HI(tie_high_T6Y26), .LO(tie_low_T6Y26));
  sky130_fd_sc_hd__conb_1 conb_T6Y27 (.HI(tie_high_T6Y27), .LO(tie_low_T6Y27));
  sky130_fd_sc_hd__conb_1 conb_T6Y28 (.HI(tie_high_T6Y28), .LO(tie_low_T6Y28));
  sky130_fd_sc_hd__conb_1 conb_T6Y29 (.HI(tie_high_T6Y29), .LO(tie_low_T6Y29));
  sky130_fd_sc_hd__conb_1 conb_T6Y3 (.HI(tie_high_T6Y3), .LO(tie_low_T6Y3));
  sky130_fd_sc_hd__conb_1 conb_T6Y30 (.HI(tie_high_T6Y30), .LO(tie_low_T6Y30));
  sky130_fd_sc_hd__conb_1 conb_T6Y31 (.HI(tie_high_T6Y31), .LO(tie_low_T6Y31));
  sky130_fd_sc_hd__conb_1 conb_T6Y32 (.HI(tie_high_T6Y32), .LO(tie_low_T6Y32));
  sky130_fd_sc_hd__conb_1 conb_T6Y33 (.HI(tie_high_T6Y33), .LO(tie_low_T6Y33));
  sky130_fd_sc_hd__conb_1 conb_T6Y34 (.HI(tie_high_T6Y34), .LO(tie_low_T6Y34));
  sky130_fd_sc_hd__conb_1 conb_T6Y35 (.HI(tie_high_T6Y35), .LO(tie_low_T6Y35));
  sky130_fd_sc_hd__conb_1 conb_T6Y36 (.HI(tie_high_T6Y36), .LO(tie_low_T6Y36));
  sky130_fd_sc_hd__conb_1 conb_T6Y37 (.HI(tie_high_T6Y37), .LO(tie_low_T6Y37));
  sky130_fd_sc_hd__conb_1 conb_T6Y38 (.HI(tie_high_T6Y38), .LO(tie_low_T6Y38));
  sky130_fd_sc_hd__conb_1 conb_T6Y39 (.HI(tie_high_T6Y39), .LO(tie_low_T6Y39));
  sky130_fd_sc_hd__conb_1 conb_T6Y4 (.HI(tie_high_T6Y4), .LO(tie_low_T6Y4));
  sky130_fd_sc_hd__conb_1 conb_T6Y40 (.HI(tie_high_T6Y40), .LO(tie_low_T6Y40));
  sky130_fd_sc_hd__conb_1 conb_T6Y41 (.HI(tie_high_T6Y41), .LO(tie_low_T6Y41));
  sky130_fd_sc_hd__conb_1 conb_T6Y42 (.HI(tie_high_T6Y42), .LO(tie_low_T6Y42));
  sky130_fd_sc_hd__conb_1 conb_T6Y43 (.HI(tie_high_T6Y43), .LO(tie_low_T6Y43));
  sky130_fd_sc_hd__conb_1 conb_T6Y44 (.HI(tie_high_T6Y44), .LO(tie_low_T6Y44));
  sky130_fd_sc_hd__conb_1 conb_T6Y45 (.HI(tie_high_T6Y45), .LO(tie_low_T6Y45));
  sky130_fd_sc_hd__conb_1 conb_T6Y46 (.HI(tie_high_T6Y46), .LO(tie_low_T6Y46));
  sky130_fd_sc_hd__conb_1 conb_T6Y47 (.HI(tie_high_T6Y47), .LO(tie_low_T6Y47));
  sky130_fd_sc_hd__conb_1 conb_T6Y48 (.HI(tie_high_T6Y48), .LO(tie_low_T6Y48));
  sky130_fd_sc_hd__conb_1 conb_T6Y49 (.HI(tie_high_T6Y49), .LO(tie_low_T6Y49));
  sky130_fd_sc_hd__conb_1 conb_T6Y5 (.HI(tie_high_T6Y5), .LO(tie_low_T6Y5));
  sky130_fd_sc_hd__conb_1 conb_T6Y50 (.HI(tie_high_T6Y50), .LO(tie_low_T6Y50));
  sky130_fd_sc_hd__conb_1 conb_T6Y51 (.HI(tie_high_T6Y51), .LO(tie_low_T6Y51));
  sky130_fd_sc_hd__conb_1 conb_T6Y52 (.HI(tie_high_T6Y52), .LO(tie_low_T6Y52));
  sky130_fd_sc_hd__conb_1 conb_T6Y53 (.HI(tie_high_T6Y53), .LO(tie_low_T6Y53));
  sky130_fd_sc_hd__conb_1 conb_T6Y54 (.HI(tie_high_T6Y54), .LO(tie_low_T6Y54));
  sky130_fd_sc_hd__conb_1 conb_T6Y55 (.HI(tie_high_T6Y55), .LO(tie_low_T6Y55));
  sky130_fd_sc_hd__conb_1 conb_T6Y56 (.HI(tie_high_T6Y56), .LO(tie_low_T6Y56));
  sky130_fd_sc_hd__conb_1 conb_T6Y57 (.HI(tie_high_T6Y57), .LO(tie_low_T6Y57));
  sky130_fd_sc_hd__conb_1 conb_T6Y58 (.HI(tie_high_T6Y58), .LO(tie_low_T6Y58));
  sky130_fd_sc_hd__conb_1 conb_T6Y59 (.HI(tie_high_T6Y59), .LO(tie_low_T6Y59));
  sky130_fd_sc_hd__conb_1 conb_T6Y6 (.HI(tie_high_T6Y6), .LO(tie_low_T6Y6));
  sky130_fd_sc_hd__conb_1 conb_T6Y60 (.HI(tie_high_T6Y60), .LO(tie_low_T6Y60));
  sky130_fd_sc_hd__conb_1 conb_T6Y61 (.HI(tie_high_T6Y61), .LO(tie_low_T6Y61));
  sky130_fd_sc_hd__conb_1 conb_T6Y62 (.HI(tie_high_T6Y62), .LO(tie_low_T6Y62));
  sky130_fd_sc_hd__conb_1 conb_T6Y63 (.HI(tie_high_T6Y63), .LO(tie_low_T6Y63));
  sky130_fd_sc_hd__conb_1 conb_T6Y64 (.HI(tie_high_T6Y64), .LO(tie_low_T6Y64));
  sky130_fd_sc_hd__conb_1 conb_T6Y65 (.HI(tie_high_T6Y65), .LO(tie_low_T6Y65));
  sky130_fd_sc_hd__conb_1 conb_T6Y66 (.HI(tie_high_T6Y66), .LO(tie_low_T6Y66));
  sky130_fd_sc_hd__conb_1 conb_T6Y67 (.HI(tie_high_T6Y67), .LO(tie_low_T6Y67));
  sky130_fd_sc_hd__conb_1 conb_T6Y68 (.HI(tie_high_T6Y68), .LO(tie_low_T6Y68));
  sky130_fd_sc_hd__conb_1 conb_T6Y69 (.HI(tie_high_T6Y69), .LO(tie_low_T6Y69));
  sky130_fd_sc_hd__conb_1 conb_T6Y7 (.HI(tie_high_T6Y7), .LO(tie_low_T6Y7));
  sky130_fd_sc_hd__conb_1 conb_T6Y70 (.HI(tie_high_T6Y70), .LO(tie_low_T6Y70));
  sky130_fd_sc_hd__conb_1 conb_T6Y71 (.HI(tie_high_T6Y71), .LO(tie_low_T6Y71));
  sky130_fd_sc_hd__conb_1 conb_T6Y72 (.HI(tie_high_T6Y72), .LO(tie_low_T6Y72));
  sky130_fd_sc_hd__conb_1 conb_T6Y73 (.HI(tie_high_T6Y73), .LO(tie_low_T6Y73));
  sky130_fd_sc_hd__conb_1 conb_T6Y74 (.HI(tie_high_T6Y74), .LO(tie_low_T6Y74));
  sky130_fd_sc_hd__conb_1 conb_T6Y75 (.HI(tie_high_T6Y75), .LO(tie_low_T6Y75));
  sky130_fd_sc_hd__conb_1 conb_T6Y76 (.HI(tie_high_T6Y76), .LO(tie_low_T6Y76));
  sky130_fd_sc_hd__conb_1 conb_T6Y77 (.HI(tie_high_T6Y77), .LO(tie_low_T6Y77));
  sky130_fd_sc_hd__conb_1 conb_T6Y78 (.HI(tie_high_T6Y78), .LO(tie_low_T6Y78));
  sky130_fd_sc_hd__conb_1 conb_T6Y79 (.HI(tie_high_T6Y79), .LO(tie_low_T6Y79));
  sky130_fd_sc_hd__conb_1 conb_T6Y8 (.HI(tie_high_T6Y8), .LO(tie_low_T6Y8));
  sky130_fd_sc_hd__conb_1 conb_T6Y80 (.HI(tie_high_T6Y80), .LO(tie_low_T6Y80));
  sky130_fd_sc_hd__conb_1 conb_T6Y81 (.HI(tie_high_T6Y81), .LO(tie_low_T6Y81));
  sky130_fd_sc_hd__conb_1 conb_T6Y82 (.HI(tie_high_T6Y82), .LO(tie_low_T6Y82));
  sky130_fd_sc_hd__conb_1 conb_T6Y83 (.HI(tie_high_T6Y83), .LO(tie_low_T6Y83));
  sky130_fd_sc_hd__conb_1 conb_T6Y84 (.HI(tie_high_T6Y84), .LO(tie_low_T6Y84));
  sky130_fd_sc_hd__conb_1 conb_T6Y85 (.HI(tie_high_T6Y85), .LO(tie_low_T6Y85));
  sky130_fd_sc_hd__conb_1 conb_T6Y86 (.HI(tie_high_T6Y86), .LO(tie_low_T6Y86));
  sky130_fd_sc_hd__conb_1 conb_T6Y87 (.HI(tie_high_T6Y87), .LO(tie_low_T6Y87));
  sky130_fd_sc_hd__conb_1 conb_T6Y88 (.HI(tie_high_T6Y88), .LO(tie_low_T6Y88));
  sky130_fd_sc_hd__conb_1 conb_T6Y89 (.HI(tie_high_T6Y89), .LO(tie_low_T6Y89));
  sky130_fd_sc_hd__conb_1 conb_T6Y9 (.HI(tie_high_T6Y9), .LO(tie_low_T6Y9));
  sky130_fd_sc_hd__conb_1 conb_T7Y0 (.HI(tie_high_T7Y0), .LO(tie_low_T7Y0));
  sky130_fd_sc_hd__conb_1 conb_T7Y1 (.HI(tie_high_T7Y1), .LO(tie_low_T7Y1));
  sky130_fd_sc_hd__conb_1 conb_T7Y10 (.HI(tie_high_T7Y10), .LO(tie_low_T7Y10));
  sky130_fd_sc_hd__conb_1 conb_T7Y11 (.HI(tie_high_T7Y11), .LO(tie_low_T7Y11));
  sky130_fd_sc_hd__conb_1 conb_T7Y12 (.HI(tie_high_T7Y12), .LO(tie_low_T7Y12));
  sky130_fd_sc_hd__conb_1 conb_T7Y13 (.HI(tie_high_T7Y13), .LO(tie_low_T7Y13));
  sky130_fd_sc_hd__conb_1 conb_T7Y14 (.HI(tie_high_T7Y14), .LO(tie_low_T7Y14));
  sky130_fd_sc_hd__conb_1 conb_T7Y15 (.HI(tie_high_T7Y15), .LO(tie_low_T7Y15));
  sky130_fd_sc_hd__conb_1 conb_T7Y16 (.HI(tie_high_T7Y16), .LO(tie_low_T7Y16));
  sky130_fd_sc_hd__conb_1 conb_T7Y17 (.HI(tie_high_T7Y17), .LO(tie_low_T7Y17));
  sky130_fd_sc_hd__conb_1 conb_T7Y18 (.HI(tie_high_T7Y18), .LO(tie_low_T7Y18));
  sky130_fd_sc_hd__conb_1 conb_T7Y19 (.HI(tie_high_T7Y19), .LO(tie_low_T7Y19));
  sky130_fd_sc_hd__conb_1 conb_T7Y2 (.HI(tie_high_T7Y2), .LO(tie_low_T7Y2));
  sky130_fd_sc_hd__conb_1 conb_T7Y20 (.HI(tie_high_T7Y20), .LO(tie_low_T7Y20));
  sky130_fd_sc_hd__conb_1 conb_T7Y21 (.HI(tie_high_T7Y21), .LO(tie_low_T7Y21));
  sky130_fd_sc_hd__conb_1 conb_T7Y22 (.HI(tie_high_T7Y22), .LO(tie_low_T7Y22));
  sky130_fd_sc_hd__conb_1 conb_T7Y23 (.HI(tie_high_T7Y23), .LO(tie_low_T7Y23));
  sky130_fd_sc_hd__conb_1 conb_T7Y24 (.HI(tie_high_T7Y24), .LO(tie_low_T7Y24));
  sky130_fd_sc_hd__conb_1 conb_T7Y25 (.HI(tie_high_T7Y25), .LO(tie_low_T7Y25));
  sky130_fd_sc_hd__conb_1 conb_T7Y26 (.HI(tie_high_T7Y26), .LO(tie_low_T7Y26));
  sky130_fd_sc_hd__conb_1 conb_T7Y27 (.HI(tie_high_T7Y27), .LO(tie_low_T7Y27));
  sky130_fd_sc_hd__conb_1 conb_T7Y28 (.HI(tie_high_T7Y28), .LO(tie_low_T7Y28));
  sky130_fd_sc_hd__conb_1 conb_T7Y29 (.HI(tie_high_T7Y29), .LO(tie_low_T7Y29));
  sky130_fd_sc_hd__conb_1 conb_T7Y3 (.HI(tie_high_T7Y3), .LO(tie_low_T7Y3));
  sky130_fd_sc_hd__conb_1 conb_T7Y30 (.HI(tie_high_T7Y30), .LO(tie_low_T7Y30));
  sky130_fd_sc_hd__conb_1 conb_T7Y31 (.HI(tie_high_T7Y31), .LO(tie_low_T7Y31));
  sky130_fd_sc_hd__conb_1 conb_T7Y32 (.HI(tie_high_T7Y32), .LO(tie_low_T7Y32));
  sky130_fd_sc_hd__conb_1 conb_T7Y33 (.HI(tie_high_T7Y33), .LO(tie_low_T7Y33));
  sky130_fd_sc_hd__conb_1 conb_T7Y34 (.HI(tie_high_T7Y34), .LO(tie_low_T7Y34));
  sky130_fd_sc_hd__conb_1 conb_T7Y35 (.HI(tie_high_T7Y35), .LO(tie_low_T7Y35));
  sky130_fd_sc_hd__conb_1 conb_T7Y36 (.HI(tie_high_T7Y36), .LO(tie_low_T7Y36));
  sky130_fd_sc_hd__conb_1 conb_T7Y37 (.HI(tie_high_T7Y37), .LO(tie_low_T7Y37));
  sky130_fd_sc_hd__conb_1 conb_T7Y38 (.HI(tie_high_T7Y38), .LO(tie_low_T7Y38));
  sky130_fd_sc_hd__conb_1 conb_T7Y39 (.HI(tie_high_T7Y39), .LO(tie_low_T7Y39));
  sky130_fd_sc_hd__conb_1 conb_T7Y4 (.HI(tie_high_T7Y4), .LO(tie_low_T7Y4));
  sky130_fd_sc_hd__conb_1 conb_T7Y40 (.HI(tie_high_T7Y40), .LO(tie_low_T7Y40));
  sky130_fd_sc_hd__conb_1 conb_T7Y41 (.HI(tie_high_T7Y41), .LO(tie_low_T7Y41));
  sky130_fd_sc_hd__conb_1 conb_T7Y42 (.HI(tie_high_T7Y42), .LO(tie_low_T7Y42));
  sky130_fd_sc_hd__conb_1 conb_T7Y43 (.HI(tie_high_T7Y43), .LO(tie_low_T7Y43));
  sky130_fd_sc_hd__conb_1 conb_T7Y44 (.HI(tie_high_T7Y44), .LO(tie_low_T7Y44));
  sky130_fd_sc_hd__conb_1 conb_T7Y45 (.HI(tie_high_T7Y45), .LO(tie_low_T7Y45));
  sky130_fd_sc_hd__conb_1 conb_T7Y46 (.HI(tie_high_T7Y46), .LO(tie_low_T7Y46));
  sky130_fd_sc_hd__conb_1 conb_T7Y47 (.HI(tie_high_T7Y47), .LO(tie_low_T7Y47));
  sky130_fd_sc_hd__conb_1 conb_T7Y48 (.HI(tie_high_T7Y48), .LO(tie_low_T7Y48));
  sky130_fd_sc_hd__conb_1 conb_T7Y49 (.HI(tie_high_T7Y49), .LO(tie_low_T7Y49));
  sky130_fd_sc_hd__conb_1 conb_T7Y5 (.HI(tie_high_T7Y5), .LO(tie_low_T7Y5));
  sky130_fd_sc_hd__conb_1 conb_T7Y50 (.HI(tie_high_T7Y50), .LO(tie_low_T7Y50));
  sky130_fd_sc_hd__conb_1 conb_T7Y51 (.HI(tie_high_T7Y51), .LO(tie_low_T7Y51));
  sky130_fd_sc_hd__conb_1 conb_T7Y52 (.HI(tie_high_T7Y52), .LO(tie_low_T7Y52));
  sky130_fd_sc_hd__conb_1 conb_T7Y53 (.HI(tie_high_T7Y53), .LO(tie_low_T7Y53));
  sky130_fd_sc_hd__conb_1 conb_T7Y54 (.HI(tie_high_T7Y54), .LO(tie_low_T7Y54));
  sky130_fd_sc_hd__conb_1 conb_T7Y55 (.HI(tie_high_T7Y55), .LO(tie_low_T7Y55));
  sky130_fd_sc_hd__conb_1 conb_T7Y56 (.HI(tie_high_T7Y56), .LO(tie_low_T7Y56));
  sky130_fd_sc_hd__conb_1 conb_T7Y57 (.HI(tie_high_T7Y57), .LO(tie_low_T7Y57));
  sky130_fd_sc_hd__conb_1 conb_T7Y58 (.HI(tie_high_T7Y58), .LO(tie_low_T7Y58));
  sky130_fd_sc_hd__conb_1 conb_T7Y59 (.HI(tie_high_T7Y59), .LO(tie_low_T7Y59));
  sky130_fd_sc_hd__conb_1 conb_T7Y6 (.HI(tie_high_T7Y6), .LO(tie_low_T7Y6));
  sky130_fd_sc_hd__conb_1 conb_T7Y60 (.HI(tie_high_T7Y60), .LO(tie_low_T7Y60));
  sky130_fd_sc_hd__conb_1 conb_T7Y61 (.HI(tie_high_T7Y61), .LO(tie_low_T7Y61));
  sky130_fd_sc_hd__conb_1 conb_T7Y62 (.HI(tie_high_T7Y62), .LO(tie_low_T7Y62));
  sky130_fd_sc_hd__conb_1 conb_T7Y63 (.HI(tie_high_T7Y63), .LO(tie_low_T7Y63));
  sky130_fd_sc_hd__conb_1 conb_T7Y64 (.HI(tie_high_T7Y64), .LO(tie_low_T7Y64));
  sky130_fd_sc_hd__conb_1 conb_T7Y65 (.HI(tie_high_T7Y65), .LO(tie_low_T7Y65));
  sky130_fd_sc_hd__conb_1 conb_T7Y66 (.HI(tie_high_T7Y66), .LO(tie_low_T7Y66));
  sky130_fd_sc_hd__conb_1 conb_T7Y67 (.HI(tie_high_T7Y67), .LO(tie_low_T7Y67));
  sky130_fd_sc_hd__conb_1 conb_T7Y68 (.HI(tie_high_T7Y68), .LO(tie_low_T7Y68));
  sky130_fd_sc_hd__conb_1 conb_T7Y69 (.HI(tie_high_T7Y69), .LO(tie_low_T7Y69));
  sky130_fd_sc_hd__conb_1 conb_T7Y7 (.HI(tie_high_T7Y7), .LO(tie_low_T7Y7));
  sky130_fd_sc_hd__conb_1 conb_T7Y70 (.HI(tie_high_T7Y70), .LO(tie_low_T7Y70));
  sky130_fd_sc_hd__conb_1 conb_T7Y71 (.HI(tie_high_T7Y71), .LO(tie_low_T7Y71));
  sky130_fd_sc_hd__conb_1 conb_T7Y72 (.HI(tie_high_T7Y72), .LO(tie_low_T7Y72));
  sky130_fd_sc_hd__conb_1 conb_T7Y73 (.HI(tie_high_T7Y73), .LO(tie_low_T7Y73));
  sky130_fd_sc_hd__conb_1 conb_T7Y74 (.HI(tie_high_T7Y74), .LO(tie_low_T7Y74));
  sky130_fd_sc_hd__conb_1 conb_T7Y75 (.HI(tie_high_T7Y75), .LO(tie_low_T7Y75));
  sky130_fd_sc_hd__conb_1 conb_T7Y76 (.HI(tie_high_T7Y76), .LO(tie_low_T7Y76));
  sky130_fd_sc_hd__conb_1 conb_T7Y77 (.HI(tie_high_T7Y77), .LO(tie_low_T7Y77));
  sky130_fd_sc_hd__conb_1 conb_T7Y78 (.HI(tie_high_T7Y78), .LO(tie_low_T7Y78));
  sky130_fd_sc_hd__conb_1 conb_T7Y79 (.HI(tie_high_T7Y79), .LO(tie_low_T7Y79));
  sky130_fd_sc_hd__conb_1 conb_T7Y8 (.HI(tie_high_T7Y8), .LO(tie_low_T7Y8));
  sky130_fd_sc_hd__conb_1 conb_T7Y80 (.HI(tie_high_T7Y80), .LO(tie_low_T7Y80));
  sky130_fd_sc_hd__conb_1 conb_T7Y81 (.HI(tie_high_T7Y81), .LO(tie_low_T7Y81));
  sky130_fd_sc_hd__conb_1 conb_T7Y82 (.HI(tie_high_T7Y82), .LO(tie_low_T7Y82));
  sky130_fd_sc_hd__conb_1 conb_T7Y83 (.HI(tie_high_T7Y83), .LO(tie_low_T7Y83));
  sky130_fd_sc_hd__conb_1 conb_T7Y84 (.HI(tie_high_T7Y84), .LO(tie_low_T7Y84));
  sky130_fd_sc_hd__conb_1 conb_T7Y85 (.HI(tie_high_T7Y85), .LO(tie_low_T7Y85));
  sky130_fd_sc_hd__conb_1 conb_T7Y86 (.HI(tie_high_T7Y86), .LO(tie_low_T7Y86));
  sky130_fd_sc_hd__conb_1 conb_T7Y87 (.HI(tie_high_T7Y87), .LO(tie_low_T7Y87));
  sky130_fd_sc_hd__conb_1 conb_T7Y88 (.HI(tie_high_T7Y88), .LO(tie_low_T7Y88));
  sky130_fd_sc_hd__conb_1 conb_T7Y89 (.HI(tie_high_T7Y89), .LO(tie_low_T7Y89));
  sky130_fd_sc_hd__conb_1 conb_T7Y9 (.HI(tie_high_T7Y9), .LO(tie_low_T7Y9));
  sky130_fd_sc_hd__conb_1 conb_T8Y0 (.HI(tie_high_T8Y0), .LO(tie_low_T8Y0));
  sky130_fd_sc_hd__conb_1 conb_T8Y1 (.HI(tie_high_T8Y1), .LO(tie_low_T8Y1));
  sky130_fd_sc_hd__conb_1 conb_T8Y10 (.HI(tie_high_T8Y10), .LO(tie_low_T8Y10));
  sky130_fd_sc_hd__conb_1 conb_T8Y11 (.HI(tie_high_T8Y11), .LO(tie_low_T8Y11));
  sky130_fd_sc_hd__conb_1 conb_T8Y12 (.HI(tie_high_T8Y12), .LO(tie_low_T8Y12));
  sky130_fd_sc_hd__conb_1 conb_T8Y13 (.HI(tie_high_T8Y13), .LO(tie_low_T8Y13));
  sky130_fd_sc_hd__conb_1 conb_T8Y14 (.HI(tie_high_T8Y14), .LO(tie_low_T8Y14));
  sky130_fd_sc_hd__conb_1 conb_T8Y15 (.HI(tie_high_T8Y15), .LO(tie_low_T8Y15));
  sky130_fd_sc_hd__conb_1 conb_T8Y16 (.HI(tie_high_T8Y16), .LO(tie_low_T8Y16));
  sky130_fd_sc_hd__conb_1 conb_T8Y17 (.HI(tie_high_T8Y17), .LO(tie_low_T8Y17));
  sky130_fd_sc_hd__conb_1 conb_T8Y18 (.HI(tie_high_T8Y18), .LO(tie_low_T8Y18));
  sky130_fd_sc_hd__conb_1 conb_T8Y19 (.HI(tie_high_T8Y19), .LO(tie_low_T8Y19));
  sky130_fd_sc_hd__conb_1 conb_T8Y2 (.HI(tie_high_T8Y2), .LO(tie_low_T8Y2));
  sky130_fd_sc_hd__conb_1 conb_T8Y20 (.HI(tie_high_T8Y20), .LO(tie_low_T8Y20));
  sky130_fd_sc_hd__conb_1 conb_T8Y21 (.HI(tie_high_T8Y21), .LO(tie_low_T8Y21));
  sky130_fd_sc_hd__conb_1 conb_T8Y22 (.HI(tie_high_T8Y22), .LO(tie_low_T8Y22));
  sky130_fd_sc_hd__conb_1 conb_T8Y23 (.HI(tie_high_T8Y23), .LO(tie_low_T8Y23));
  sky130_fd_sc_hd__conb_1 conb_T8Y24 (.HI(tie_high_T8Y24), .LO(tie_low_T8Y24));
  sky130_fd_sc_hd__conb_1 conb_T8Y25 (.HI(tie_high_T8Y25), .LO(tie_low_T8Y25));
  sky130_fd_sc_hd__conb_1 conb_T8Y26 (.HI(tie_high_T8Y26), .LO(tie_low_T8Y26));
  sky130_fd_sc_hd__conb_1 conb_T8Y27 (.HI(tie_high_T8Y27), .LO(tie_low_T8Y27));
  sky130_fd_sc_hd__conb_1 conb_T8Y28 (.HI(tie_high_T8Y28), .LO(tie_low_T8Y28));
  sky130_fd_sc_hd__conb_1 conb_T8Y29 (.HI(tie_high_T8Y29), .LO(tie_low_T8Y29));
  sky130_fd_sc_hd__conb_1 conb_T8Y3 (.HI(tie_high_T8Y3), .LO(tie_low_T8Y3));
  sky130_fd_sc_hd__conb_1 conb_T8Y30 (.HI(tie_high_T8Y30), .LO(tie_low_T8Y30));
  sky130_fd_sc_hd__conb_1 conb_T8Y31 (.HI(tie_high_T8Y31), .LO(tie_low_T8Y31));
  sky130_fd_sc_hd__conb_1 conb_T8Y32 (.HI(tie_high_T8Y32), .LO(tie_low_T8Y32));
  sky130_fd_sc_hd__conb_1 conb_T8Y33 (.HI(tie_high_T8Y33), .LO(tie_low_T8Y33));
  sky130_fd_sc_hd__conb_1 conb_T8Y34 (.HI(tie_high_T8Y34), .LO(tie_low_T8Y34));
  sky130_fd_sc_hd__conb_1 conb_T8Y35 (.HI(tie_high_T8Y35), .LO(tie_low_T8Y35));
  sky130_fd_sc_hd__conb_1 conb_T8Y36 (.HI(tie_high_T8Y36), .LO(tie_low_T8Y36));
  sky130_fd_sc_hd__conb_1 conb_T8Y37 (.HI(tie_high_T8Y37), .LO(tie_low_T8Y37));
  sky130_fd_sc_hd__conb_1 conb_T8Y38 (.HI(tie_high_T8Y38), .LO(tie_low_T8Y38));
  sky130_fd_sc_hd__conb_1 conb_T8Y39 (.HI(tie_high_T8Y39), .LO(tie_low_T8Y39));
  sky130_fd_sc_hd__conb_1 conb_T8Y4 (.HI(tie_high_T8Y4), .LO(tie_low_T8Y4));
  sky130_fd_sc_hd__conb_1 conb_T8Y40 (.HI(tie_high_T8Y40), .LO(tie_low_T8Y40));
  sky130_fd_sc_hd__conb_1 conb_T8Y41 (.HI(tie_high_T8Y41), .LO(tie_low_T8Y41));
  sky130_fd_sc_hd__conb_1 conb_T8Y42 (.HI(tie_high_T8Y42), .LO(tie_low_T8Y42));
  sky130_fd_sc_hd__conb_1 conb_T8Y43 (.HI(tie_high_T8Y43), .LO(tie_low_T8Y43));
  sky130_fd_sc_hd__conb_1 conb_T8Y44 (.HI(tie_high_T8Y44), .LO(tie_low_T8Y44));
  sky130_fd_sc_hd__conb_1 conb_T8Y45 (.HI(tie_high_T8Y45), .LO(tie_low_T8Y45));
  sky130_fd_sc_hd__conb_1 conb_T8Y46 (.HI(tie_high_T8Y46), .LO(tie_low_T8Y46));
  sky130_fd_sc_hd__conb_1 conb_T8Y47 (.HI(tie_high_T8Y47), .LO(tie_low_T8Y47));
  sky130_fd_sc_hd__conb_1 conb_T8Y48 (.HI(tie_high_T8Y48), .LO(tie_low_T8Y48));
  sky130_fd_sc_hd__conb_1 conb_T8Y49 (.HI(tie_high_T8Y49), .LO(tie_low_T8Y49));
  sky130_fd_sc_hd__conb_1 conb_T8Y5 (.HI(tie_high_T8Y5), .LO(tie_low_T8Y5));
  sky130_fd_sc_hd__conb_1 conb_T8Y50 (.HI(tie_high_T8Y50), .LO(tie_low_T8Y50));
  sky130_fd_sc_hd__conb_1 conb_T8Y51 (.HI(tie_high_T8Y51), .LO(tie_low_T8Y51));
  sky130_fd_sc_hd__conb_1 conb_T8Y52 (.HI(tie_high_T8Y52), .LO(tie_low_T8Y52));
  sky130_fd_sc_hd__conb_1 conb_T8Y53 (.HI(tie_high_T8Y53), .LO(tie_low_T8Y53));
  sky130_fd_sc_hd__conb_1 conb_T8Y54 (.HI(tie_high_T8Y54), .LO(tie_low_T8Y54));
  sky130_fd_sc_hd__conb_1 conb_T8Y55 (.HI(tie_high_T8Y55), .LO(tie_low_T8Y55));
  sky130_fd_sc_hd__conb_1 conb_T8Y56 (.HI(tie_high_T8Y56), .LO(tie_low_T8Y56));
  sky130_fd_sc_hd__conb_1 conb_T8Y57 (.HI(tie_high_T8Y57), .LO(tie_low_T8Y57));
  sky130_fd_sc_hd__conb_1 conb_T8Y58 (.HI(tie_high_T8Y58), .LO(tie_low_T8Y58));
  sky130_fd_sc_hd__conb_1 conb_T8Y59 (.HI(tie_high_T8Y59), .LO(tie_low_T8Y59));
  sky130_fd_sc_hd__conb_1 conb_T8Y6 (.HI(tie_high_T8Y6), .LO(tie_low_T8Y6));
  sky130_fd_sc_hd__conb_1 conb_T8Y60 (.HI(tie_high_T8Y60), .LO(tie_low_T8Y60));
  sky130_fd_sc_hd__conb_1 conb_T8Y61 (.HI(tie_high_T8Y61), .LO(tie_low_T8Y61));
  sky130_fd_sc_hd__conb_1 conb_T8Y62 (.HI(tie_high_T8Y62), .LO(tie_low_T8Y62));
  sky130_fd_sc_hd__conb_1 conb_T8Y63 (.HI(tie_high_T8Y63), .LO(tie_low_T8Y63));
  sky130_fd_sc_hd__conb_1 conb_T8Y64 (.HI(tie_high_T8Y64), .LO(tie_low_T8Y64));
  sky130_fd_sc_hd__conb_1 conb_T8Y65 (.HI(tie_high_T8Y65), .LO(tie_low_T8Y65));
  sky130_fd_sc_hd__conb_1 conb_T8Y66 (.HI(tie_high_T8Y66), .LO(tie_low_T8Y66));
  sky130_fd_sc_hd__conb_1 conb_T8Y67 (.HI(tie_high_T8Y67), .LO(tie_low_T8Y67));
  sky130_fd_sc_hd__conb_1 conb_T8Y68 (.HI(tie_high_T8Y68), .LO(tie_low_T8Y68));
  sky130_fd_sc_hd__conb_1 conb_T8Y69 (.HI(tie_high_T8Y69), .LO(tie_low_T8Y69));
  sky130_fd_sc_hd__conb_1 conb_T8Y7 (.HI(tie_high_T8Y7), .LO(tie_low_T8Y7));
  sky130_fd_sc_hd__conb_1 conb_T8Y70 (.HI(tie_high_T8Y70), .LO(tie_low_T8Y70));
  sky130_fd_sc_hd__conb_1 conb_T8Y71 (.HI(tie_high_T8Y71), .LO(tie_low_T8Y71));
  sky130_fd_sc_hd__conb_1 conb_T8Y72 (.HI(tie_high_T8Y72), .LO(tie_low_T8Y72));
  sky130_fd_sc_hd__conb_1 conb_T8Y73 (.HI(tie_high_T8Y73), .LO(tie_low_T8Y73));
  sky130_fd_sc_hd__conb_1 conb_T8Y74 (.HI(tie_high_T8Y74), .LO(tie_low_T8Y74));
  sky130_fd_sc_hd__conb_1 conb_T8Y75 (.HI(tie_high_T8Y75), .LO(tie_low_T8Y75));
  sky130_fd_sc_hd__conb_1 conb_T8Y76 (.HI(tie_high_T8Y76), .LO(tie_low_T8Y76));
  sky130_fd_sc_hd__conb_1 conb_T8Y77 (.HI(tie_high_T8Y77), .LO(tie_low_T8Y77));
  sky130_fd_sc_hd__conb_1 conb_T8Y78 (.HI(tie_high_T8Y78), .LO(tie_low_T8Y78));
  sky130_fd_sc_hd__conb_1 conb_T8Y79 (.HI(tie_high_T8Y79), .LO(tie_low_T8Y79));
  sky130_fd_sc_hd__conb_1 conb_T8Y8 (.HI(tie_high_T8Y8), .LO(tie_low_T8Y8));
  sky130_fd_sc_hd__conb_1 conb_T8Y80 (.HI(tie_high_T8Y80), .LO(tie_low_T8Y80));
  sky130_fd_sc_hd__conb_1 conb_T8Y81 (.HI(tie_high_T8Y81), .LO(tie_low_T8Y81));
  sky130_fd_sc_hd__conb_1 conb_T8Y82 (.HI(tie_high_T8Y82), .LO(tie_low_T8Y82));
  sky130_fd_sc_hd__conb_1 conb_T8Y83 (.HI(tie_high_T8Y83), .LO(tie_low_T8Y83));
  sky130_fd_sc_hd__conb_1 conb_T8Y84 (.HI(tie_high_T8Y84), .LO(tie_low_T8Y84));
  sky130_fd_sc_hd__conb_1 conb_T8Y85 (.HI(tie_high_T8Y85), .LO(tie_low_T8Y85));
  sky130_fd_sc_hd__conb_1 conb_T8Y86 (.HI(tie_high_T8Y86), .LO(tie_low_T8Y86));
  sky130_fd_sc_hd__conb_1 conb_T8Y87 (.HI(tie_high_T8Y87), .LO(tie_low_T8Y87));
  sky130_fd_sc_hd__conb_1 conb_T8Y88 (.HI(tie_high_T8Y88), .LO(tie_low_T8Y88));
  sky130_fd_sc_hd__conb_1 conb_T8Y89 (.HI(tie_high_T8Y89), .LO(tie_low_T8Y89));
  sky130_fd_sc_hd__conb_1 conb_T8Y9 (.HI(tie_high_T8Y9), .LO(tie_low_T8Y9));
  sky130_fd_sc_hd__conb_1 conb_T9Y0 (.HI(tie_high_T9Y0), .LO(tie_low_T9Y0));
  sky130_fd_sc_hd__conb_1 conb_T9Y1 (.HI(tie_high_T9Y1), .LO(tie_low_T9Y1));
  sky130_fd_sc_hd__conb_1 conb_T9Y10 (.HI(tie_high_T9Y10), .LO(tie_low_T9Y10));
  sky130_fd_sc_hd__conb_1 conb_T9Y11 (.HI(tie_high_T9Y11), .LO(tie_low_T9Y11));
  sky130_fd_sc_hd__conb_1 conb_T9Y12 (.HI(tie_high_T9Y12), .LO(tie_low_T9Y12));
  sky130_fd_sc_hd__conb_1 conb_T9Y13 (.HI(tie_high_T9Y13), .LO(tie_low_T9Y13));
  sky130_fd_sc_hd__conb_1 conb_T9Y14 (.HI(tie_high_T9Y14), .LO(tie_low_T9Y14));
  sky130_fd_sc_hd__conb_1 conb_T9Y15 (.HI(tie_high_T9Y15), .LO(tie_low_T9Y15));
  sky130_fd_sc_hd__conb_1 conb_T9Y16 (.HI(tie_high_T9Y16), .LO(tie_low_T9Y16));
  sky130_fd_sc_hd__conb_1 conb_T9Y17 (.HI(tie_high_T9Y17), .LO(tie_low_T9Y17));
  sky130_fd_sc_hd__conb_1 conb_T9Y18 (.HI(tie_high_T9Y18), .LO(tie_low_T9Y18));
  sky130_fd_sc_hd__conb_1 conb_T9Y19 (.HI(tie_high_T9Y19), .LO(tie_low_T9Y19));
  sky130_fd_sc_hd__conb_1 conb_T9Y2 (.HI(tie_high_T9Y2), .LO(tie_low_T9Y2));
  sky130_fd_sc_hd__conb_1 conb_T9Y20 (.HI(tie_high_T9Y20), .LO(tie_low_T9Y20));
  sky130_fd_sc_hd__conb_1 conb_T9Y21 (.HI(tie_high_T9Y21), .LO(tie_low_T9Y21));
  sky130_fd_sc_hd__conb_1 conb_T9Y22 (.HI(tie_high_T9Y22), .LO(tie_low_T9Y22));
  sky130_fd_sc_hd__conb_1 conb_T9Y23 (.HI(tie_high_T9Y23), .LO(tie_low_T9Y23));
  sky130_fd_sc_hd__conb_1 conb_T9Y24 (.HI(tie_high_T9Y24), .LO(tie_low_T9Y24));
  sky130_fd_sc_hd__conb_1 conb_T9Y25 (.HI(tie_high_T9Y25), .LO(tie_low_T9Y25));
  sky130_fd_sc_hd__conb_1 conb_T9Y26 (.HI(tie_high_T9Y26), .LO(tie_low_T9Y26));
  sky130_fd_sc_hd__conb_1 conb_T9Y27 (.HI(tie_high_T9Y27), .LO(tie_low_T9Y27));
  sky130_fd_sc_hd__conb_1 conb_T9Y28 (.HI(tie_high_T9Y28), .LO(tie_low_T9Y28));
  sky130_fd_sc_hd__conb_1 conb_T9Y29 (.HI(tie_high_T9Y29), .LO(tie_low_T9Y29));
  sky130_fd_sc_hd__conb_1 conb_T9Y3 (.HI(tie_high_T9Y3), .LO(tie_low_T9Y3));
  sky130_fd_sc_hd__conb_1 conb_T9Y30 (.HI(tie_high_T9Y30), .LO(tie_low_T9Y30));
  sky130_fd_sc_hd__conb_1 conb_T9Y31 (.HI(tie_high_T9Y31), .LO(tie_low_T9Y31));
  sky130_fd_sc_hd__conb_1 conb_T9Y32 (.HI(tie_high_T9Y32), .LO(tie_low_T9Y32));
  sky130_fd_sc_hd__conb_1 conb_T9Y33 (.HI(tie_high_T9Y33), .LO(tie_low_T9Y33));
  sky130_fd_sc_hd__conb_1 conb_T9Y34 (.HI(tie_high_T9Y34), .LO(tie_low_T9Y34));
  sky130_fd_sc_hd__conb_1 conb_T9Y35 (.HI(tie_high_T9Y35), .LO(tie_low_T9Y35));
  sky130_fd_sc_hd__conb_1 conb_T9Y36 (.HI(tie_high_T9Y36), .LO(tie_low_T9Y36));
  sky130_fd_sc_hd__conb_1 conb_T9Y37 (.HI(tie_high_T9Y37), .LO(tie_low_T9Y37));
  sky130_fd_sc_hd__conb_1 conb_T9Y38 (.HI(tie_high_T9Y38), .LO(tie_low_T9Y38));
  sky130_fd_sc_hd__conb_1 conb_T9Y39 (.HI(tie_high_T9Y39), .LO(tie_low_T9Y39));
  sky130_fd_sc_hd__conb_1 conb_T9Y4 (.HI(tie_high_T9Y4), .LO(tie_low_T9Y4));
  sky130_fd_sc_hd__conb_1 conb_T9Y40 (.HI(tie_high_T9Y40), .LO(tie_low_T9Y40));
  sky130_fd_sc_hd__conb_1 conb_T9Y41 (.HI(tie_high_T9Y41), .LO(tie_low_T9Y41));
  sky130_fd_sc_hd__conb_1 conb_T9Y42 (.HI(tie_high_T9Y42), .LO(tie_low_T9Y42));
  sky130_fd_sc_hd__conb_1 conb_T9Y43 (.HI(tie_high_T9Y43), .LO(tie_low_T9Y43));
  sky130_fd_sc_hd__conb_1 conb_T9Y44 (.HI(tie_high_T9Y44), .LO(tie_low_T9Y44));
  sky130_fd_sc_hd__conb_1 conb_T9Y45 (.HI(tie_high_T9Y45), .LO(tie_low_T9Y45));
  sky130_fd_sc_hd__conb_1 conb_T9Y46 (.HI(tie_high_T9Y46), .LO(tie_low_T9Y46));
  sky130_fd_sc_hd__conb_1 conb_T9Y47 (.HI(tie_high_T9Y47), .LO(tie_low_T9Y47));
  sky130_fd_sc_hd__conb_1 conb_T9Y48 (.HI(tie_high_T9Y48), .LO(tie_low_T9Y48));
  sky130_fd_sc_hd__conb_1 conb_T9Y49 (.HI(tie_high_T9Y49), .LO(tie_low_T9Y49));
  sky130_fd_sc_hd__conb_1 conb_T9Y5 (.HI(tie_high_T9Y5), .LO(tie_low_T9Y5));
  sky130_fd_sc_hd__conb_1 conb_T9Y50 (.HI(tie_high_T9Y50), .LO(tie_low_T9Y50));
  sky130_fd_sc_hd__conb_1 conb_T9Y51 (.HI(tie_high_T9Y51), .LO(tie_low_T9Y51));
  sky130_fd_sc_hd__conb_1 conb_T9Y52 (.HI(tie_high_T9Y52), .LO(tie_low_T9Y52));
  sky130_fd_sc_hd__conb_1 conb_T9Y53 (.HI(tie_high_T9Y53), .LO(tie_low_T9Y53));
  sky130_fd_sc_hd__conb_1 conb_T9Y54 (.HI(tie_high_T9Y54), .LO(tie_low_T9Y54));
  sky130_fd_sc_hd__conb_1 conb_T9Y55 (.HI(tie_high_T9Y55), .LO(tie_low_T9Y55));
  sky130_fd_sc_hd__conb_1 conb_T9Y56 (.HI(tie_high_T9Y56), .LO(tie_low_T9Y56));
  sky130_fd_sc_hd__conb_1 conb_T9Y57 (.HI(tie_high_T9Y57), .LO(tie_low_T9Y57));
  sky130_fd_sc_hd__conb_1 conb_T9Y58 (.HI(tie_high_T9Y58), .LO(tie_low_T9Y58));
  sky130_fd_sc_hd__conb_1 conb_T9Y59 (.HI(tie_high_T9Y59), .LO(tie_low_T9Y59));
  sky130_fd_sc_hd__conb_1 conb_T9Y6 (.HI(tie_high_T9Y6), .LO(tie_low_T9Y6));
  sky130_fd_sc_hd__conb_1 conb_T9Y60 (.HI(tie_high_T9Y60), .LO(tie_low_T9Y60));
  sky130_fd_sc_hd__conb_1 conb_T9Y61 (.HI(tie_high_T9Y61), .LO(tie_low_T9Y61));
  sky130_fd_sc_hd__conb_1 conb_T9Y62 (.HI(tie_high_T9Y62), .LO(tie_low_T9Y62));
  sky130_fd_sc_hd__conb_1 conb_T9Y63 (.HI(tie_high_T9Y63), .LO(tie_low_T9Y63));
  sky130_fd_sc_hd__conb_1 conb_T9Y64 (.HI(tie_high_T9Y64), .LO(tie_low_T9Y64));
  sky130_fd_sc_hd__conb_1 conb_T9Y65 (.HI(tie_high_T9Y65), .LO(tie_low_T9Y65));
  sky130_fd_sc_hd__conb_1 conb_T9Y66 (.HI(tie_high_T9Y66), .LO(tie_low_T9Y66));
  sky130_fd_sc_hd__conb_1 conb_T9Y67 (.HI(tie_high_T9Y67), .LO(tie_low_T9Y67));
  sky130_fd_sc_hd__conb_1 conb_T9Y68 (.HI(tie_high_T9Y68), .LO(tie_low_T9Y68));
  sky130_fd_sc_hd__conb_1 conb_T9Y69 (.HI(tie_high_T9Y69), .LO(tie_low_T9Y69));
  sky130_fd_sc_hd__conb_1 conb_T9Y7 (.HI(tie_high_T9Y7), .LO(tie_low_T9Y7));
  sky130_fd_sc_hd__conb_1 conb_T9Y70 (.HI(tie_high_T9Y70), .LO(tie_low_T9Y70));
  sky130_fd_sc_hd__conb_1 conb_T9Y71 (.HI(tie_high_T9Y71), .LO(tie_low_T9Y71));
  sky130_fd_sc_hd__conb_1 conb_T9Y72 (.HI(tie_high_T9Y72), .LO(tie_low_T9Y72));
  sky130_fd_sc_hd__conb_1 conb_T9Y73 (.HI(tie_high_T9Y73), .LO(tie_low_T9Y73));
  sky130_fd_sc_hd__conb_1 conb_T9Y74 (.HI(tie_high_T9Y74), .LO(tie_low_T9Y74));
  sky130_fd_sc_hd__conb_1 conb_T9Y75 (.HI(tie_high_T9Y75), .LO(tie_low_T9Y75));
  sky130_fd_sc_hd__conb_1 conb_T9Y76 (.HI(tie_high_T9Y76), .LO(tie_low_T9Y76));
  sky130_fd_sc_hd__conb_1 conb_T9Y77 (.HI(tie_high_T9Y77), .LO(tie_low_T9Y77));
  sky130_fd_sc_hd__conb_1 conb_T9Y78 (.HI(tie_high_T9Y78), .LO(tie_low_T9Y78));
  sky130_fd_sc_hd__conb_1 conb_T9Y79 (.HI(tie_high_T9Y79), .LO(tie_low_T9Y79));
  sky130_fd_sc_hd__conb_1 conb_T9Y8 (.HI(tie_high_T9Y8), .LO(tie_low_T9Y8));
  sky130_fd_sc_hd__conb_1 conb_T9Y80 (.HI(tie_high_T9Y80), .LO(tie_low_T9Y80));
  sky130_fd_sc_hd__conb_1 conb_T9Y81 (.HI(tie_high_T9Y81), .LO(tie_low_T9Y81));
  sky130_fd_sc_hd__conb_1 conb_T9Y82 (.HI(tie_high_T9Y82), .LO(tie_low_T9Y82));
  sky130_fd_sc_hd__conb_1 conb_T9Y83 (.HI(tie_high_T9Y83), .LO(tie_low_T9Y83));
  sky130_fd_sc_hd__conb_1 conb_T9Y84 (.HI(tie_high_T9Y84), .LO(tie_low_T9Y84));
  sky130_fd_sc_hd__conb_1 conb_T9Y85 (.HI(tie_high_T9Y85), .LO(tie_low_T9Y85));
  sky130_fd_sc_hd__conb_1 conb_T9Y86 (.HI(tie_high_T9Y86), .LO(tie_low_T9Y86));
  sky130_fd_sc_hd__conb_1 conb_T9Y87 (.HI(tie_high_T9Y87), .LO(tie_low_T9Y87));
  sky130_fd_sc_hd__conb_1 conb_T9Y88 (.HI(tie_high_T9Y88), .LO(tie_low_T9Y88));
  sky130_fd_sc_hd__conb_1 conb_T9Y89 (.HI(tie_high_T9Y89), .LO(tie_low_T9Y89));
  sky130_fd_sc_hd__conb_1 conb_T9Y9 (.HI(tie_high_T9Y9), .LO(tie_low_T9Y9));
  sky130_fd_sc_hd__clkinv_4 cts_buf_0 (.A(clk_cts_root), .X(clk_cts_n0));
  sky130_fd_sc_hd__clkinv_4 cts_buf_1 (.A(clk_cts_root), .X(clk_cts_n1));
  sky130_fd_sc_hd__clkinv_4 cts_buf_10 (.A(clk_cts_root), .X(clk_cts_n10));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_11 (.A(clk_cts_root), .X(clk_cts_n11));
  sky130_fd_sc_hd__clkinv_4 cts_buf_12 (.A(clk_cts_root), .X(clk_cts_n12));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_13 (.A(clk_cts_root), .X(clk_cts_n13));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_14 (.A(clk_cts_root), .X(clk_cts_n14));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_15 (.A(clk_cts_root), .X(clk_cts_n15));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_16 (.A(clk_cts_root), .X(clk_cts_n16));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_17 (.A(clk_cts_root), .X(clk_cts_n17));
  sky130_fd_sc_hd__clkinv_4 cts_buf_18 (.A(clk_cts_root), .X(clk_cts_n18));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_19 (.A(clk_cts_root), .X(clk_cts_n19));
  sky130_fd_sc_hd__clkinv_4 cts_buf_2 (.A(clk_cts_root), .X(clk_cts_n2));
  sky130_fd_sc_hd__clkinv_4 cts_buf_20 (.A(clk_cts_root), .X(clk_cts_n20));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_21 (.A(clk_cts_root), .X(clk_cts_n21));
  sky130_fd_sc_hd__clkinv_4 cts_buf_22 (.A(clk_cts_root), .X(clk_cts_n22));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_23 (.A(clk_cts_root), .X(clk_cts_n23));
  sky130_fd_sc_hd__clkinv_4 cts_buf_24 (.A(clk_cts_root), .X(clk_cts_n24));
  sky130_fd_sc_hd__clkinv_4 cts_buf_25 (.A(clk_cts_root), .X(clk_cts_n25));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_26 (.A(clk_cts_root), .X(clk_cts_n26));
  sky130_fd_sc_hd__clkinv_4 cts_buf_27 (.A(clk_cts_root), .X(clk_cts_n27));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_28 (.A(clk_cts_root), .X(clk_cts_n28));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_29 (.A(clk_cts_root), .X(clk_cts_n29));
  sky130_fd_sc_hd__clkinv_4 cts_buf_3 (.A(clk_cts_root), .X(clk_cts_n3));
  sky130_fd_sc_hd__clkinv_4 cts_buf_4 (.A(clk_cts_root), .X(clk_cts_n4));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_5 (.A(clk_cts_root), .X(clk_cts_n5));
  sky130_fd_sc_hd__clkinv_4 cts_buf_6 (.A(clk_cts_root), .X(clk_cts_n6));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_7 (.A(clk_cts_root), .X(clk_cts_n7));
  sky130_fd_sc_hd__clkbuf_4 cts_buf_8 (.A(clk_cts_root), .X(clk_cts_n8));
  sky130_fd_sc_hd__clkinv_4 cts_buf_9 (.A(clk_cts_root), .X(clk_cts_n9));

endmodule
